
`timescale 1ns/1ns
module u_jp2k_9(
    flush_over, zero_plane_number, codeblock_counter, 
    wr_clk, rd_clk, rst, rst_syn, data_from_mq, 
    cal_truncation_point_start, compression_ratio, 
    pass_plane, word_last_flag_plane_sp, 
    word_last_flag_plane_mp, word_last_flag_plane_cp, 
    one_codeblock_over, pass_error_plane_sp, 
    pass_error_plane_mp, pass_error_plane_cp, 


    target_slope, codeblock_shift_over, cal_truncation_point_over, 
    output_to_ram, buffer_all_over, 
    lram_write_en, lram_address_wr, target_byte_number
);

	parameter aDkQEysUQMjSKApaeshi=14,
		WORD_WIDTH=18;


	input flush_over;
	input [3:0]zero_plane_number;
	input [7:0]codeblock_counter;
	input wr_clk;
	input rd_clk;
	input rst;
	input rst_syn;
	input [15:0]data_from_mq;
	input cal_truncation_point_start;
	
	input [2:0]compression_ratio;
	input [1:0]pass_plane;
	input word_last_flag_plane_sp;
	input word_last_flag_plane_mp;
	input word_last_flag_plane_cp;
	input one_codeblock_over;
	input [30:0]pass_error_plane_sp;
	input [30:0]pass_error_plane_mp;
	input [30:0]pass_error_plane_cp;



	output [8:0]target_slope;
	output codeblock_shift_over;
	output cal_truncation_point_over;
	output [WORD_WIDTH-1:0]output_to_ram;
	output buffer_all_over;
	output lram_write_en;
	output [aDkQEysUQMjSKApaeshi-1:0]lram_address_wr;
	output [19:0]target_byte_number;

	wire TLXWChymSkORZZFunpRb;
	wire FuMFDshlwPAZNriIzdKA;
	wire codeblock_shift_over;
	wire ytSqxoZpMDkNRuAUbZDc;
	wire [1:0]nhadPSkgCafxNJCdwkKp;
	wire cal_truncation_point_over;
	wire jMCVmjFKEszeMFGJPhDT;
	wire [37:0]CxvpyAhqMqQXTLpXgdOB;
	wire [37:0]JBFuaKfGSzMztOCsXGjt;
	wire [15:0]iGrqtIPPBFPUhGunhSdw;
    wire [15:0]CZceBwenUmhgWecdrVuw;
    wire [15:0]FODhltaveISdQIJPBJhJ;
    wire [15:0]mBUfUweOiYOTkxaNfvqZ;
    wire [15:0]XCEBnusbPkduEdkiHxFK;
    wire [15:0]UKLUuuVquDsMMMMhkoJV;
	wire	[7:0]	LkKGICfCcYyYLBJKtucQ; 
	wire	[7:0]	SupobFuabxSWuLFQTEEe; 
	wire	[7:0]	BUOYkUPXSUGjGnnMOiLz; 
	wire	[7:0]	tOmHmkYobOhcasHrvveC; 
	wire	[7:0]	HMRNTVVBwfsQwiaIOdeu; 
	wire	[7:0]	hGCZylpOryFfZNhxLZOH; 
	wire GVEVAzxUWjnkLWGcHbCC;
	wire artgRMUHHAMMXysfVQxf;
	wire ZOkiujEkXjtpgkcONTax;
	wire CcBPKbMCVTPpuzcHaNNl;
	wire QcQmUnoklSTURFcjjsxj;
	wire MQgLtHVUbOxalviVAmNV;
	wire qUkWgSUxlHDGwaShnpJD;
    wire AKnQHFnRxMsayGvtbpFT;
    wire EdvpzeTpOWEloDTnpLTm;
    wire vWFpyuXCRPPETqWnXLgO;
    wire dbsLvjpjMhdBsPiUgbjQ;
    wire oXZLEogkFzslyJXIZmAm;
	wire [38:0]rczbRGCFDOHKNTiwObwc;
	wire [38:0]OHenhlDjGfxNrcoKTDTe;
	wire [7:0]FssIYlUsXIkosBplffKR;
	wire [7:0]fvbJniljSNczcXeDYDTv;
	wire [2:0]uoqQSqkDyZwtvuETruXA;
	wire [2:0]AnaDOfYtVBlpyqvNRuwL;
	wire [2:0]irdAYQxVjzyKmWopQQGP;


	reg [5:0]daVvNjfwJBQRozThYCld;
	reg [3:0]XtrJUtwJnzBPPMzRDosc;
	reg buffer_all_over;
	reg nQAnZVgoKyprBQAdRCfA;
	reg wEtGDzRjafclnvKxgCSP;
	reg [2:0]YfuArrGnpBUyrJxEvVgI;
	reg [3:0]tQSdMsmQOoDjgNvoiCmq;
	reg LrLbKGgLtBSEzbICsDNb;
	reg DnfnMYzlPFszZtXlGDhW;
	reg NhvFLRUduFzxNErEsMee;
	reg FGUJmfBLDaAxYUKmfnyF;
	reg [8:0]target_slope;
	reg [8:0]qgkpXRmlTwkWNutDGWMM;
	reg [19:0]GVfnzKKftzXfxeBqPQMD;
	reg [19:0]target_byte_number;
	reg lram_write_en;
	reg [aDkQEysUQMjSKApaeshi-1:0]lram_address_wr;
	reg XmWQfEltjOUqcNLDCtfd;
	reg pyhAjCtAJLKGgXMclzgY;
	reg MPFTDVkljwqlROSuxXcP;
	reg [29:0]ESEFEoPuTgYdvrsaqlOz;
	reg [4:0]ARQLJGuTZBnFJHXDoAkT;
	reg [4:0]gStNdqadtalDMswfRuqW;                         
	reg [4:0]euqWRDzuVBfSvNZlbygs;                     
	reg [5:0]XWSDWJpZwWFziLcqAlai;
	reg [7:0]CHmFHLXDhsSOMWPfgbXw;
	reg eojmGbYrZBcDvhuhplcn;
	reg [17:0]output_to_ram;
	reg [7:0]qaVKoOckmCbhBtxSbviM;
	reg [7:0]wKozjyqvbxpraCSNGCJY;
	reg [8:0]OhIQvlSNredlAvEzVwlD;
	reg [8:0]bVNTszDvPimBrKwNycBW;
	reg [7:0]CTJvELJpTGwHTCgirGVs;
	reg [15:0]aSItvOfWsSQOkHOHMzuM;
	reg [29:0]oEDxWLutHlOkrCgasnsy;
	reg kAXRTBBnwMdFccjIlXSw;

	
	reg [29:0]RdPhRZcalGKJvMOvrAIh;
	reg [29:0]xMPttPagqqqJUKztQdOZ;
	reg [29:0]YCteCIAKCruidjpeILHG;
	reg [29:0]nxlEkFPUCwQVbIQJmgbx;
	reg [29:0]SVzsQtfHGQqXqNoloxvo;
	reg [29:0]vMLEZaXExwsFFvafFmfc;
	reg [3:0]MNhKBwmQfBNRRoCGsGYL  ;//{{{
	reg [3:0]CZUlnpSgUmTCmXxNawKq  ;
	reg [3:0]GCKDpTZdSkziHIHQTHTY  ;
	reg [3:0]TbggffYtMBhiLSACnOtm  ;
	reg [3:0]QMFreKPqLMtYHbzgqBQA  ;
	reg [3:0]NlcVQzrrHSpHBCrquBjt  ;
	reg [3:0]FSYqURbHbEaesQcTkdrx  ;
	reg [3:0]qEtkygphCMCbDqrWtklY  ;
	reg [3:0]TLjaqwEsoHtrvWTBQRsK  ;
	reg [3:0]cYsREsbuuQNtJwVuIQtc ;
	reg [3:0]IADijSHmLDuBqTQJOxSa ;
	reg [3:0]BhAYLsocIYeStsZZVTUF ;
	reg [3:0]WQWSkTgEaMFMXPEsFHwg ;
	reg [3:0]WVikipTMfwFUtPMyACXK ;
	reg [3:0]dXrKEPxqSBOppMxaytbW ;
	reg [3:0]NnjJwuwNoVWroSgcnSsE ;
	reg [3:0]ASCWICejFoBbZHMJMVyD ;
	reg [3:0]twyoccXqjNTyiiCHZKgQ ;
	reg [3:0]xvRCARkQSEXoZFEiGfjC ;
	reg [3:0]JjLGddxBYbYmoYBVjdju ;
	reg [3:0]xyvvBnpUfpnejSAdOrIU ;
	reg [3:0]LNWqJGCGvJkqDqnyFdST ;
	reg [3:0]XXnujvRmwKtqZZbYXNom ;
	reg [3:0]rdgcYAhdMEGqsgkVVhHB ;
	reg [3:0]bcCzAdPYbGFOdbqFGtNY ;
	reg [3:0]MRTHuncHaQWNXrTdnjLu ;
	reg [3:0]ZqxWPnvGQEisPGNSDkWt ;
	reg [3:0]jLboxjBIZGftrbnYaDHz ;
	reg [3:0]XPHrltKlkTYeddIYErlL ;
	reg [3:0]DwnEuDbYEGceHCFfntWU ;
	reg [3:0]AhXRxsizDLdrPCSJbgvu ;
	reg [3:0]dRLKJNMhCWjmYIXyBBMS ;
	reg [3:0]qKakmPsWXvxWDjopwmhd ;
	reg [3:0]OfKBQrlHgohHRFQMqPuX ;
	reg [3:0]OMUVfbzXJtBmpgGUlWIN ;
	reg [3:0]pRjKNldSGgrOVpMtRdhl ;
	reg [3:0]FzItXojZYuRrQPYroXqa ;
	reg [3:0]tiASKMApdODRGubKCrIk ;
	reg [3:0]AofWIQWGCHGeAWxyBSnX ;
	reg [3:0]BVZJHRZIRDJUNzlhOXNj ;
	reg [3:0]MJngMbRNrQAqZKOoJbfA ;
	reg [3:0]LKEbaiUcnUkcdhTlxIWn ;
	reg [3:0]PIdKWDjIZqdVETXVKUyz ;
	reg [3:0]TeweoifYlvYAXegPEOev ;
	reg [3:0]aHdPRBehEsBXhVSVEVGI ;
	reg [3:0]EHDzFoGEUiKMcpmeZndO ;
	reg [3:0]iGWdFxfLkcoPAfSnTRiW ;
	reg [3:0]OgwvxakMlGIDTjsTTTrF ;
	reg [3:0]hweOwCSFFCFpnLABsNDz ;
	reg [3:0]kFILldZgHWqtwHcEyrEz ;
	reg [8:0]BHxWpRKaPloRmedcGnVS ;
	reg [8:0]jEDhTzjvJVSeQkYxJusx ;
	reg [8:0]nVWwCingLJiAmNkXNBse ;
	reg [8:0]hdQpCNCsCpWxWjyDHYIf ;
	reg [8:0]mYfjBwhqQaPjGDGuVzVT ;
	reg [8:0]sPdTjZhZROmcYPkfxnHK ;
	reg [8:0]VOSkkJBkJQjLTSFCXXZG ;
	reg [8:0]wnDMhVWFcihAknOuJWgt ;
	reg [8:0]ZJYNMlOSJujZtBMVfIcG ;
	reg [8:0]cUQgUjrarAoCxWvadhrh ;
	reg [8:0]ayPBmMeTERtfSkylBBkl ;
	reg [8:0]zjiIArXGbkjgPxxXfPxg ;
	reg [8:0]YERHnxdykgyyioNNZJSQ ;
	reg [8:0]rNuBwbgCniYGlSgOMCnE ;
	reg [8:0]VjtVxkxLZrdVPkMsyEqe ;
	reg [8:0]fFwIafFNLTVTiIeJUZOi ;
	reg [8:0]JofSpHHAILpRCvnGOmzf ;
	reg [8:0]OeYMhMfjeDdvkecHiLUT ;
	reg [8:0]tVOTCptQSOpsjFBXiksw ;
	reg [8:0]AhXuWEaSPuUvIcwDuFWr ;
	reg [8:0]ekQuaIqPJyasZNSLaQOo ;
	reg [8:0]osvtoSWcIuWcmvZruLsS ;
	reg [8:0]BzXYfwLRzqKLxtfxvmZC ;
	reg [8:0]tgVDzxwqtPquEcvdvFrC ;
	reg [8:0]DzNsyDbNrzFrSyvQMHnd ;
	reg [8:0]iOnjZhBOoaDLaXXeVrwx ;
	reg [8:0]XwvNGtBVJXErWQRUuqBI ;
	reg [8:0]JJgTPGsdUTcAdufkeJgK ;
	reg [8:0]TfnRFMUqcGKfwYVkrOcp ;
	reg [8:0]kuHTqKTEGHJGjcgKEkCF ;
	reg [8:0]FfvTBiXNEwWARzrRMUYh ;
	reg [8:0]VMfdRrsDolDymeMDbscN ;
	reg [8:0]iPuXoTiWLBGZVYAHGaYO ;
	reg [8:0]BaxkmTikPlEanrOALJQn ;
	reg [8:0]TGPYgdsEOqsHqlpqyhVp ;
	reg [8:0]VZaWDekOPjcbcuLkmTCK ;
	reg [8:0]ceSSpUnFGIqusvzAQYyv ;
	reg [8:0]KkgZHqKRoBphLNurbXZv ;
	reg [8:0]BVfKHJmimWhfvhFZYdJC ;
	reg [8:0]XWIoNGOmiUqZuWDNerJA ;
	reg [8:0]ymZNoaOSvkuMNFrKCZJc ;
	reg [8:0]JtPboWbpZfxqTBEEDYyf ;
	reg [8:0]NIzOkTmOrsmtdJpYgwkn ;
	reg [8:0]HPBVjcjYzqThfAZsuBko ;
	reg [8:0]RtOUSNvLjifycdHERnsH ;
	reg [8:0]RHqjRVMUmlsTYhhiTxqt ;
	reg [8:0]irQWRPjnSymTgyEWfOeV ;
	reg [8:0]gHMMxJFDpgQtSoSKsfzc ;
	reg [8:0]XrXzzUeQwqtdbHighLXh ;
	reg [8:0]VXesUOJyNaYiksaASUmr; 
	reg [8:0]MjDYzSbWZYtgtBPeFxFX; 
	reg [8:0]QocIghyhzPXBoGjaFxEW; 
	reg [8:0]aNNRDAQndlQbuwTNoeBC; 
	reg [8:0]ganwYnOuHsVFGlnGQGGf; 
	reg [8:0]TmUIbPULspEIyexiGCHU; 
	reg [8:0]GrWFHsoruHLBTofZiNlc; 
	reg [8:0]HemnvXRItkGWOQQBARSS; 
	reg [8:0]crDvxwhExTyEkehZAJBR; 
	reg [8:0]vqFRiEdZYIvaYIjwIZPo; 
	reg [8:0]RiyBtzLqNImqdjYXxYLF; 
	reg [8:0]QAZelRxmduKrKymXyprg; 
	reg [8:0]IixlIEeyecDFQCcIcXFK; 
	reg [8:0]CahtEzYLkeeOsdRKBvoI; 
	reg [8:0]hXvwCaJPKLmTlGnIqShO; 
	reg [8:0]ZapMeflJnJGQFrDdnzZx; 
	reg [8:0]tEZVPsZbWePhmBDkYbkW; 
	reg [8:0]VKIhSekuVtyFcvuoBpZH; 
	reg [8:0]HHissIgZPvjjCfGzZWgP; 
	reg [8:0]ZthEdVQnyODdQJpzqpDX; 
	reg [8:0]ZvVAYFyMKYuJjjuLlssM; 
	reg [8:0]BDVfxjBZqdgfpcXaqSxS; 
	reg [8:0]SYPrSAmIZhepjzRpfAbW; 
	reg [8:0]bheecNbLIfuKFYksBrvM; 
	reg [8:0]LoFfmBmHEBmQlYvRihJx; 
	reg [8:0]RAqkMVQdcCkZqHQrYhTY; 
	reg [8:0]JwazcQrhGdLokRSxMIPy; 
	reg [8:0]NHwKTvStgXGxecepjZCb; 
	reg [8:0]iFhOAEkrfnWgTHHMCrAr; 
	reg [8:0]KoZvZIhKhWDYlgwhYWfH; 
	reg [8:0]xqkVQlUmzixmBBOWsogM; 
	reg [8:0]mZcXpTwcGpwcsXaAXzJZ; 
	reg [8:0]tBkJHywSnDHjCloeCKQN; 
	reg [8:0]rtIOwgMybhKPbMtTkPHH; 
	reg [8:0]ULvOWCBpLiqodnUiPZne; 
	reg [8:0]UeCtXzcgpZHmscgLWNgU; 
	reg [8:0]NchYslfTwDoJDaIhKQld; 
	reg [8:0]vdLrgmXBDTPmGWwCZgJK; 
	reg [8:0]fypmfZbmWDbDCXEismjU; 
	reg [8:0]FEgAuSjALENQXZOiGFUZ; 
	reg [8:0]hUaTrhFAshrngFoHaXaJ; 
	reg [8:0]avmhenqBbGIfSBAIabaF; 
	reg [8:0]IlmCWYrxdJVqIQywKmAF; 
	reg [8:0]GXKZdRvGRyUFWKyHVAFD; 
	reg [8:0]PExEfPxznaZHuROUSmfc; 
	reg [8:0]DoWtmJCIdGMmwEInsyhi; 
	reg [8:0]AtkWXjDVDEZLaumbWZzI; 
	reg [8:0]HvOvrGAvaPTzYsRxiQFa; 
	reg [8:0]rwPuhbqaLGfEsTZJaDhF; 
	reg [8:0]YphfuswJNWiAbvgWEfjm; 
	reg [8:0]YhTJCIYfjiXccwQDAncB; 
	reg [8:0]KaDxyGuuayhqIxIwbGQG; 
	reg [8:0]SCcERabQMmiRZhSuKFqS; 
	reg [8:0]ASVDnraQDtLQhInOEyVK; 
	reg [8:0]RzDedJWchbeEickgtFOM; 
	reg [8:0]qBWQIFhDbnPbANWZJPUR; 
	reg [8:0]ONSywhEkLUpjhsBVzOEr; 
	reg [8:0]SiWXyZwStCTfnlFxLPQx; 
	reg [8:0]ljlzMOdncFtIKCHtOsVQ; 
	reg [8:0]sBtkXBZAHFHDVqMZHZdd; 
	reg [8:0]ZNywgghYzvszBznGurzE; 
	reg [8:0]giByCXZhzRJrKpUfJiYx; 
	reg [8:0]NOzoIRcSVgyFREyzzHqs; 
	reg [8:0]hvcttLppSPcVixtVRHqN; 
	reg [8:0]NXURaWZymtMESRzASoml; 
	reg [8:0]OGJwXjhBDuVzMrVxGthI; 
	reg [8:0]tDHSWWPwhDHPIdkjEtEW; 
	reg [8:0]spPgPLHCbVgdzOmJFakw; 
	reg [8:0]NCLfdSDEGhGvIWQaIuMS; 
	reg [8:0]NfdfbTCtNjYFDeLLecMe; 
	reg [8:0]xIHGyzqgFJSHmjAJEkTk; 
	reg [8:0]ffdnbvLvbNGfaiXRKcYD; 
	reg [8:0]dDkKlvBKHVNSwGZicnzg; 
	reg [8:0]sTYRbAXFBXVNlExKcFRO; 
	reg [8:0]QYcegkQFzbKFzvlPxGeR; 
	reg [8:0]WCbGOTtDaZUdMPlupDBN; 
	reg [8:0]kNoeoxFOMGDTBbVzHlLM; 
	reg [8:0]pcsafTpJQiyaKivHSiiO; 
	reg [8:0]HhgKJaIdyWwhlApPzTKC; 
	reg [8:0]LgxgHDHmFYbeGgXVWgvC; 
	reg [8:0]cKBOWdNoOXhznBHdAwlu; 
	reg [8:0]KASZraJCWhbAUtfwnLfk; 
	reg [8:0]AGPbOkqoDAYNiAUBxYWb; 
	reg [8:0]QePGiiHhRVKoAUkzEcSD; 
	reg [8:0]ULkqQHcjawmJPPtzcPCS; 
	reg [8:0]gVMkJmsMEYFtEfiuwaKj; 
	reg [8:0]yHFGaozymIVZZMqtzLDd; 
	reg [8:0]XyhfMHNDiNoQgejMGALx; 
	reg [8:0]zWhpxSLccsmBmQBUhbQT; 
	reg [8:0]xKWgakKpWyTQyBrwYCIS; 
	reg [8:0]UkOdSdYxtcxumOakhLgx; 
	reg [8:0]nhnBLnxptnOVgbmRStCU; 
	reg [8:0]UmXpnIjWZNlfEPEYcDTn; 
	reg [8:0]deblhPqNAplcidEXSGqw; 
	reg [8:0]GgkZJHLDkhyFsCCzuqLa; 
	reg [8:0]pKDUrDrLLWTOdoUxvsyF; 
	reg [8:0]JrQYFpYwpBTANpnTvLiU; 
	reg [8:0]KencLjTnnSFqjwbVxqJg; 
	reg [8:0]TXuaPuUIuhCkLiMhEKiF; 
	reg [8:0]aAhmLslHTfVKwKSRWVtp; 
	reg [8:0]NJEYMnPHSmEVDftsqzQE; 
	reg [8:0]ByBgtRovBsKUVHUQEzwk; 
	reg [8:0]pcCSuYOgcgRTEfyKANVf; 
	reg [8:0]OOJGXLeAUSSWDwWKvqMN; 
	reg [8:0]xzObOtBnVrtyMpWImLGp; 
	reg [8:0]fPvbFzCudNRdKXFIwPTW; 
	reg [8:0]UCBlEpPTGRkqheRhrmew; 
	reg [8:0]rxGiYeZlkdsRNUfrmDKO; 
	reg [8:0]BRDRPJjxjaVvUmeEcabW; 
	reg [8:0]twevQhSVcRXlOWMZGHZH; 
	reg [8:0]hsPTsFDtcTjmyeddHGwC; 
	reg [8:0]SnXYHdlnJsKNjOCDlAdk; 
	reg [8:0]fzPjNCWXNlBXDEixcMfx; 
	reg [8:0]MzxTqhCibhKKovZUinvJ; 
	reg [8:0]UjBCIuRFDGUvCwBBwjtv; 
	reg [8:0]WLvkMHkFFjSeXeCMFLqU; 
	reg [8:0]OdXRCGgZgKmtknFfVeGS; 
	reg [8:0]YTagschVaYsVmCoZyGxw; 
	reg [8:0]uBDeqwBeWjkFnJPifZac; 
	reg [8:0]ChqdVbAPIMvlcdCLZFDM; 
	reg [8:0]xVhIWQmsjbKYhycXOZZj; 
	reg [8:0]moXSbLoysxSoGKFutzbo; 
	reg [8:0]pFrrbOJSlADGwICgxTdA; 
	reg [8:0]eFKOOLSSWbJGsojVvoDI; 
	reg [8:0]CjkyDsWsnyjeHKnTfjoz; 
	reg [8:0]ikgPtqNHSxOonFiPgvOK; 
	reg [8:0]JzYgxPBzYqfsNCHdKwWT; 
	reg [8:0]rYlFPAhuURCPKCloqLOG; 
	reg [8:0]PQEjeJZSeiJdTNkqSiiS; 
	reg [8:0]MSaMrnCOKHvvWjrvrLVh; 
	reg [8:0]bZovfeygdcHHRKfkxfHl; 
	reg [8:0]ATkQsyvByLEkPXEmCGoF; 
	reg [8:0]uBtJXFukNYPqTHWppmdv; 
	reg [8:0]soNzOmONAzHkpLFWdCtg; 
	reg [8:0]lLJeyDbtTaFvkSfqLcWK; 
	reg [8:0]lMFLPXTVXadwnVsRrAPI; 
	reg [8:0]WPsXEglrQBPoHLKokyap; 
	reg [8:0]RqjRxpMaojbkWLGINNMj; 
	reg [8:0]CcpgUvVvfmeEoXXGYlgz; 
	reg [8:0]yNeJpDTKbQScFfOFsIMP; 
	reg [8:0]uVWYpFOIjqHtdFWqJLJL; 
	reg [8:0]vCLJZIRyvOOZpamupbmS; 
	reg [8:0]JiRCGeWXVDSjvohYatoO; 
	reg [8:0]JXVeYnVHSdAGpxmDHgjf; 
	reg [8:0]iXlLoGyimBUgUkjZoGvT; 
	reg [8:0]JrBVZVJGLbQlQIuxVRMO; 
	reg [8:0]MZLrRshlRErhPsqJeccP; 
	reg [8:0]KddqRkJXVvlRHkpsKNQL; 
	reg [8:0]eKWoIeUrKiPbRIhuWEla; 
	reg [8:0]JRsyUSbxyBGBNdlJquOD; 
	reg [8:0]mobFFnIZQLEDGamGRCMQ; 
	reg [8:0]MIfRQTaujrTsVSIdukaO; 
	reg [8:0]qQxKziPkMaoHyxLiZQNv; 
	reg [8:0]SbGofGNBnFvEqTbzCMDT; 
	reg [8:0]eAyuUdQDmhsyVqUkrWtf; 
	reg [8:0]xcrfMbSpXdXRmlkuZRPx; 
	reg [8:0]BKSeIpcsVISDrrWyloru; 
	reg [8:0]cFxrUFXVhwbgFamPfIXu; 
	reg [8:0]EawSFufNSOZZHKtrbfDb; 
	reg [8:0]TtHHtKtzZHIcJuWziTSX; 
	reg [8:0]KAQFclKTjvNuQpWZONVn; 
	reg [8:0]zdDIxzPkCVYUHKycUMxS; 
	reg [8:0]yRWhBghWQtDlHOXzOKHV; 
	reg [8:0]xzEZrlRsvTQMlJcdcoBA; 
	reg [8:0]omKttYZtWwSNmJfXmNhw; 
	reg [8:0]TJsrTmKBrLuIryymjrla; 
	reg [8:0]UQIvtuLZLyNrLBcITiBh; 
	reg [8:0]dewJijMNQrULKORvfOPu; 
	reg [8:0]fFCHqQnaXGJtQcWhDHoo; 
	reg [8:0]lDVujeiDOsfmAcgTJEeH; 
	reg [8:0]tHYVLHNrDsWBBiksZJSh; 
	reg [8:0]YGcrryHhhucPWCRpoXpV; 
	reg [8:0]vhaFurczuHuVJndQizpm; 
	reg [8:0]bAUZnBUzAeFxTBCaAwBD; 
	reg [8:0]SJSSeEtWLefcHjjHknTt; 
	reg [8:0]RrXElmqzMleQDmHbRetu; 
	reg [8:0]RiwCfvabTaSgTyqQQkNP; 
	reg [8:0]ijLmWvKcGWYkfmVliDIH; 
	reg [8:0]JhZCVmRnYDVfDuTgaJBq; 
	reg [8:0]MmtedWLnvMwKkqgwBoYk; 
	reg [8:0]xNONPhZsuWCOqfHyKvVw; 
	reg [8:0]UYtsWPGzDLbsLPHFFzpM; 
	reg [8:0]HaIozTBrCuKZJRqUpAty; 
	reg [8:0]ihhBdoTzqImqsCjVxwKM; 
	reg [8:0]LPKCNZYNtyFJTUiKvFKI; 
	reg [8:0]VcDzTcOFndjUjhnRfxTN; 
	reg [8:0]ScSvdbbLcbwcpTKFudIt; 
	reg [8:0]ZFOGopcNcymIuYXsiiRw; 
	reg [8:0]zVAojGgdEwSIpPjTZZId; 
	reg [8:0]qwGWpRzKYsDLRvxcxAAH; 
	reg [8:0]WPkpODdzyINGGhuwZyoF; 
	reg [8:0]BaxiLnGgFxSKHVKkEWrL; 
	reg [8:0]cChsgcLGnvNEmegZREam; 
	reg [8:0]FRCWHcmIuMUUWgdYMzWu; 
	reg [8:0]QDYrIGBlnoXdNCUflHOP; 
	reg [8:0]zzYTnLgksIjwqZSweXMf; 
	reg [8:0]cWljGAlocPwsnrDyMjHO; 
	reg [8:0]JPYOnWGSGjFuHZfQBaEZ; 
	reg [8:0]VzfYJEwelHYPMpUSDmsC; 
	reg [8:0]XYQGKDohhXYVCeaCtmre; 
	reg [3:0]GbajCDnxXLGTStnsYsds; 
	reg [3:0]THlQvXwjkuLqdcMtPxBy; 
	reg [3:0]avkJIgYNFpvoyRkxaMTC; 
	reg [3:0]yhgnNUWIhVDlrtUDGEZn; 
	reg [3:0]lHvULbFfwhQgtqfjhwzH; 
	reg [3:0]TymwlUFeZUaLhFoWTZzU; 
	reg [3:0]obAWtmAwdFBYPXQlSuSy; 
	reg [3:0]VBJGcheVZYcxGpvcuBoi; 
	reg [3:0]NpcOSbiIpOcdgCjboENs; 
	reg [3:0]PiHYPPmDrZQNPnlqBFSt; 
	reg [3:0]rOXoAhCRFHntxISYSkye; 
	reg [3:0]IsXHeZVJKogNnFFfJwvx; 
	reg [3:0]BtfuDWbiQheMoNKySKtm; 
	reg [3:0]lsMUeaCgYLjCPUiUXaIc; 
	reg [3:0]kTdnGvNmLrhbepFdhZCh; 
	reg [3:0]vKbnovNlLRioZoJsQunL; 
	reg [3:0]nXBrtwwgIArkXUbHKAye; 
	reg [3:0]czvIYhYPaYPpRHUBJMFc; 
	reg [3:0]nsezjQWxmqwzmxCwosDv; 
	reg [3:0]ruIyZIesSthmxIaXEtrJ; 
	reg [3:0]cXQjLxPFTWRBhlJmdxUJ; 
	reg [3:0]GPoMmfciZsakCXuJMdbD; 
	reg [3:0]sZUCFycPxeatsZozmHJN; 
	reg [3:0]XbnmwpButuNSkogDlbQb; 
	reg [3:0]wdkDXnIkWnpQMmswGQeU; 
	reg [3:0]KpEHEcApUpQBvCLoAeYT; 
	reg [3:0]KsaghLmgaRvpRfCktbJZ; 
	reg [3:0]lZVGNfUlVmsuLbJxnQDA; 
	reg [3:0]rMBkqrLcKhflEMUYxGkE; 
	reg [3:0]wMlYFxkSbZTCTvhQOIei; 
	reg [3:0]WQGVbnQQZGQWVmpcxvbb; 
	reg [3:0]AzsKalhmBYUitbArLbcU; 
	reg [3:0]ekrMWzROxYoWtRpdbLZH; 
	reg [3:0]uLMmObkZiwzDlReqMwJN; 
	reg [3:0]eAEEsZkRTlfXOeEdICRO; 
	reg [3:0]DyXCiZssIzbywKGAbIwY; 
	reg [3:0]wBOVUPcFUWzhOUKDlJVa; 
	reg [3:0]BCsgCSHvysHWLteqbRMX; 
	reg [3:0]FrvVghZEElOfAJGPEURk; 
	reg [3:0]DHNpdfPdlvcIeMhPYCBD; 
	reg [3:0]ByKBiFClfZeeoBwNqVdH; 
	reg [3:0]muXlkjUrAqYazTUUGcVg; 
	reg [3:0]rZlIolWetZZffpSrlMAn; 
	reg [3:0]fCxfzzVrwjVhwiuAOpOD; 
	reg [3:0]VHDrEEGVFWccsKXzbEjD; 
	reg [3:0]pgbmZFwAnGMkExuHZexG; 
	reg [3:0]CYTIFZXRYHDOwAOpYhTY; 
	reg [3:0]hzujftnKaamrwjRBenpS; 
	reg [3:0]DwBiXGPwomcqrFUiwGKO; 
	reg [3:0]TxOTbaXnfvTWWAEMVKsT; 
	reg [3:0]VBPMSBgUzhZWqifRFXLt; 
	reg [3:0]fBEMznDkaUpJbucpUFUs; 
	reg [3:0]RXuUWWKfwotmzMaIdOHs; 
	reg [3:0]DScSrBltRCaJuMKRHxjp; 
	reg [3:0]yKhNJjIQvjuuxuKGtNvD; 
	reg [3:0]MBLbhXLxXGZHZERKIoYb; 
	reg [3:0]AiFthZhNPfZiXSnyPCOt; 
	reg [3:0]uDpYTElkHJsWMgegRIkv; 
	reg [3:0]LqJHECWMJlDdyFDTTZZH; 
	reg [3:0]ohfsyAOCKLVNdUfnlZGT; 
	reg [3:0]MOoDdDePAGBzQbLCZlwX; 
	reg [3:0]MHLazVdHgoSmGTltAxsJ; 
	reg [3:0]CYSqcBzpHDXSSATrgQjL; 
	reg [3:0]rPKZMoWgFDpDSJXXQmEU; 
	reg [3:0]hniufLGfdzmHbDIvsTIo; 
	reg [3:0]wTfPVycgpDcgGCOQhJjH; 
	reg [3:0]lcOMvsbHZmIJccXoDkqZ; 
	reg [3:0]UKirjTCurmcGUGGogrnh; 
	reg [3:0]KVLRCNcgwgdezgxdbtiz; 
	reg [3:0]ISUkQBFCDDhkmXDnEdVT; 
	reg [3:0]wLiUXxuAUdxCuAoAbUxH; 
	reg [3:0]vQNMUmgdbJJDFKzsjqLK; 
	reg [3:0]PPaVHoPQXNFqYDIgCroQ; 
	reg [3:0]fZmgOJpwMcdeRjEcecxZ; 
	reg [3:0]pXxRQDEgUJLwgwAsNvmV; 
	reg [3:0]JWyFVCrskBwarfgMzbIK; 
	reg [3:0]nLMIykvKsueQiebJRjaB; 
	reg [3:0]MwUAnLVNdEpwKFXarSrE; 
	reg [3:0]rwKFeNNlWzDutFvKudZd; 
	reg [3:0]YFTuhpacOohGrtlEUgyn; 
	reg [3:0]orsjfJIPQQvjIhvrnfZT; 
	reg [3:0]beooHOrejCcWcSXDuAMs; 
	reg [3:0]wLFqLqnhtGKyjhXVaXLu; 
	reg [3:0]VhlEwlgxfirfMpIAJZhE; 
	reg [3:0]ybSCwixJTEhXYyRpEeDj; 
	reg [3:0]PLAwknGzfcioZVaFOQCX; 
	reg [3:0]WdDdHRBJZdBPCxmYbWdk; 
	reg [3:0]BIxIzsQvWljjGYxMCQtS; 
	reg [3:0]TZYUrtPvAdyOAezlYVJO; 
	reg [3:0]qPqZhRZBobhmAXNGrsmh; 
	reg [3:0]BCGaGkllXBcyohBosHqS; 
	reg [3:0]pcgiabuotmBHXKOYDDAq; 
	reg [3:0]VidvAsXIfsppEpKtZeYc; 
	reg [3:0]lGfaCxQtDihDBzWEuyaH; 
	reg [3:0]ucwrtDfHQDZIjkmTmCvN; 
	reg [3:0]dayIzRpYaQRnEjXynbCm; 
	reg [3:0]vqgpItmCwuhiwKZyFXMt; 
	reg [3:0]FnVEwsGKlXZfUqxZGqHn; 
	reg [3:0]bitnzrgsExKEWSXnsRZq; 
	reg [3:0]eYsNwIgUOqnSppAZBKfW; 
	reg [3:0]FXTNpbkOJRifihZRkFUk; 
	reg [3:0]UCyPKegIVHgIqztViRHP; 
	reg [3:0]urwbynurHojveDuzQAqY; 
	reg [3:0]djsdiJHbeUEoOocTIVAL; 
	reg [3:0]juEeWiBDxjlSPOBoDWca; 
	reg [3:0]ZfhQiwfaJoKgwqVVBKhf; 
	reg [3:0]SNnVNrhdPUfxhixiespl; 
	reg [3:0]cHHoYqPSIzoxFEuXvNLY; 
	reg [3:0]hLpCUWbILJOjqbDhVEwn; 
	reg [3:0]itXQCyFacJzvPyzfGwVe; 
	reg [3:0]iujmIQQClXPYAKjueUBD; 
	reg [3:0]BjdcbpGuKPxnpZzFTfte; 
	reg [3:0]ZQFzyLJsVraTCGkqQcZA; 
	reg [3:0]fADZyEOwTyWvSQFgOnwG; 
	reg [3:0]xbhqvpXrDTlnyBNQeAlC; 
	reg [3:0]usigvHtlPqTHmByMEGLy; 
	reg [3:0]EqRnSoIxQaLPlCNmpBmq; 
	reg [3:0]VzsEzvUFwafgXDXiMnOI; 
	reg [3:0]qjQChEpAPSbKmoDGRppN; 
	reg [3:0]XBdmfGxuWrXGMBFOANKF; 
	reg [3:0]iHWmgCopJntOccGPObxn; 
	reg [3:0]eeoTbTyuwxPCsjuUGnLj; 
	reg [3:0]MkxrURKJtUzHVTfBwhoO; 
	reg [3:0]USFkaPtDBVOjbGpLXKUX; 
	reg [3:0]xcBSpPXNgyeMCKwBcsxX; 
	reg [3:0]APZhwjfiYOuKluWEaTIj; 
	reg [3:0]eiYeGwmYgODBCzcNuNtn; 
	reg [3:0]rmoQVcRSrSeskIibJzCc; 
	reg [3:0]AzSDmFqniQGEkrUvtcQd; 
	reg [3:0]BYQMYRDRDKXGHnLYQyKL; 
	reg [3:0]iYaojeeenaSObFkfIEyS; 
	reg [3:0]OvjWCALXGQonpSVNSUDx; 
	reg [3:0]QNSQONiKmlvpucXZsAKo; 
	reg [3:0]RKLbOFQSgMkwEdftvnBQ; 
	reg [3:0]hoPvrLDkwXFTkYESCUcp; 
	reg [3:0]hShwACbdYktXmGxyazAM; 
	reg [3:0]puehHutFkvCRvoGqbSYp; 
	reg [3:0]CSpvXCVkXjBnWvAFEiDG; 
	reg [3:0]GBnbMGmdJLNqPHpTRJqo; 
	reg [3:0]PQFlqUWXvhfFTKRniEDA; 
	reg [3:0]mNQfwTdWpUOnxIhbTYfU; 
	reg [3:0]ldQowZgtPeXlzjFcyWQl; 
	reg [3:0]HYWHYpKWyjTHzWIzGNeE; 
	reg [3:0]vsHmuANStIQsYgoNHsHw; 
	reg [3:0]tYWmIUymjXADFjUmKFpP; 
	reg [3:0]OQmggBTvOqhAXBiDJeaP; 
	reg [3:0]EFcUAERFHbivPwgHAMQa; 
	reg [3:0]jpbydIYGKyCwhjgemImi; 
	reg [3:0]OVYjPuZDVHOTTeuFPkrT; 
	reg [3:0]DqhwOfIUxBzsVSgEjWzC; 
	reg [3:0]plztNCDwyKBliboMvXKs; 
	reg [3:0]GojVETmCGfWcYwVYimBv; 
	reg [3:0]aogDiFiAXQqphSrsQbJV; 
	reg [3:0]rCOKgSoVLfXaUWFdsBnJ; 
	reg [3:0]ZuONZDcmHxALaUULMEAA; 
	reg [3:0]KIjEeYrBOSrzUMqGYBsV; 
	reg [3:0]ZBocacKljeyYorCiQgzQ; 
	reg [3:0]mqazMnBgYnlLqLRzaNYx; 
	reg [3:0]oyfKvpCwkpoCCxTglCJr; 
	reg [3:0]NGNEGckWnRLaqnjOKOmx; 
	reg [3:0]cVWqyzzrUUodYFbrorBz; 
	reg [3:0]RjwugczIYXEQzzmUrnYh; 
	reg [3:0]lEqWgKBWIbLvYwrXeDtN; 
	reg [3:0]DhnZhzYLzUMXzuxLMdpR; 
	reg [3:0]WwogGcAbNuwPRaXHfllR; 
	reg [3:0]fymbKnqnRYaHIRuPXxle; 
	reg [3:0]nJWkhXEkUmrasSyMThpL; 
	reg [3:0]qXNWBYTrrKKKGSroThrT; 
	reg [3:0]OWgmvdYcTEmvwkEuDkJS; 
	reg [3:0]urpaOisfjSiDXEZoTBsG; 
	reg [3:0]mveotDylkopgLZJFFBVl; 
	reg [3:0]CCXECvtOeIBEOFePtIRw; 
	reg [3:0]iYYwLjjGMjLikfxxrxIB; 
	reg [3:0]BJhcDugYXUoZuTXYBzJg; 
	reg [3:0]wpEZHrezpouBVvAiIOpn; 
	reg [3:0]omjfRcaEwaSdXWjgQYUv; 
	reg [3:0]aWXCrpICnOAsyXgkDTDT; 
	reg [3:0]HjXRkNnhDmrrYeoZLfga; 
	reg [3:0]zDWiKpAenkhcNZIBSNiT; 
	reg [3:0]UfyNbuBOwMXEdumKnlqN; 
	reg [9:0]LYSwVHbgNGVrAkuDLmxY; 

	



	parameter tqCfMxDxNMUeAVjaKWqL=0,
		FIND_FIRST_PASS=1,
		CAL_SLOPE_1=2,
		CAL_SLOPE_2=3,
		CAL_SLOPE_3=4,
		SHIFT_PASS_FIRST_HEADER=5,
		SHIFT_PASS_SECOND_HEADER=6,
		SHIFT_CODESTREAM=7,
		NEXT_PASS=8,
		PASS_OVER=9, 
		CAL_TRUNCATION_POINT=10,
		CAL_TRUNCATION_POINT_OVER=11,
		BUFFER=12,
		WAITING_WRITE_OVER=13,
		SHIFT_OVER_FLAG=14,
		ONE_EMPTY_CODEBLOCK_OVER=15;

	assign codeblock_shift_over=wEtGDzRjafclnvKxgCSP&&nQAnZVgoKyprBQAdRCfA||gStNdqadtalDMswfRuqW==ONE_EMPTY_CODEBLOCK_OVER;
	assign cal_truncation_point_over=(gStNdqadtalDMswfRuqW==CAL_TRUNCATION_POINT_OVER); 
	
	always@(posedge rd_clk or negedge rst)
	begin
	    if(!rst)
			target_slope<=0;
		else if(rst_syn)
			target_slope<=0;
		else if(jMCVmjFKEszeMFGJPhDT&&lram_address_wr==480)
			target_slope<=1;
		else if(ytSqxoZpMDkNRuAUbZDc)
			target_slope<=481-lram_address_wr;    
	end
	
	always@(posedge rd_clk or negedge rst)
	begin
	    if(!rst)
			lram_address_wr<=0;
		else if(rst_syn)
			lram_address_wr<=0;
		else if(buffer_all_over)  
			lram_address_wr<=0;
		else if(lram_write_en||jMCVmjFKEszeMFGJPhDT)
			lram_address_wr<=lram_address_wr+1;     
	end
	
	always@(posedge rd_clk or negedge rst)
	begin
	    if(!rst)
			output_to_ram<=0;
		else if(rst_syn)
			output_to_ram<=0;
		else 
		begin
			case(gStNdqadtalDMswfRuqW)
				SHIFT_PASS_FIRST_HEADER:output_to_ram<={2'b11,codeblock_counter,CHmFHLXDhsSOMWPfgbXw[7:0]};
				SHIFT_PASS_SECOND_HEADER:output_to_ram<={nhadPSkgCafxNJCdwkKp[1:0],tQSdMsmQOoDjgNvoiCmq[3:0],3'b0,OhIQvlSNredlAvEzVwlD[8:0]};
				SHIFT_CODESTREAM:output_to_ram<={2'b00,aSItvOfWsSQOkHOHMzuM};
				SHIFT_OVER_FLAG:output_to_ram<={2'b11,16'hffff};
			endcase
		end
	end
	

	always@(posedge rd_clk or negedge rst)
	begin
		if(!rst)
			daVvNjfwJBQRozThYCld<=0;
		else if(rst_syn)
			daVvNjfwJBQRozThYCld<=0;
		else if(nQAnZVgoKyprBQAdRCfA&&one_codeblock_over)   
			daVvNjfwJBQRozThYCld<=daVvNjfwJBQRozThYCld+1;
		else if(gStNdqadtalDMswfRuqW==ONE_EMPTY_CODEBLOCK_OVER)
			daVvNjfwJBQRozThYCld<=daVvNjfwJBQRozThYCld-1;
	end
	
	always@(posedge rd_clk or negedge rst)
	begin
		if(!rst)
			XtrJUtwJnzBPPMzRDosc<=0;
		else if(rst_syn)
			XtrJUtwJnzBPPMzRDosc<=XtrJUtwJnzBPPMzRDosc+1;
		else if(codeblock_shift_over)
			XtrJUtwJnzBPPMzRDosc<=0;
		else if(flush_over)
			XtrJUtwJnzBPPMzRDosc<=XtrJUtwJnzBPPMzRDosc+1;      
	end
	
	always@(posedge rd_clk or negedge rst)
	begin
		if(!rst)
			buffer_all_over<=0;
		else if(rst_syn)
			buffer_all_over<=0;
		else if(gStNdqadtalDMswfRuqW==SHIFT_OVER_FLAG)
			buffer_all_over<=1;
		else buffer_all_over<=0;
	end
	always@(posedge rd_clk or negedge rst)
	begin
	    if(!rst)
			YfuArrGnpBUyrJxEvVgI<=0;
		else if(rst_syn)
			YfuArrGnpBUyrJxEvVgI<=0;
		else if(YfuArrGnpBUyrJxEvVgI==5)
			YfuArrGnpBUyrJxEvVgI<=0;
		else if(gStNdqadtalDMswfRuqW==WAITING_WRITE_OVER)
			YfuArrGnpBUyrJxEvVgI<=YfuArrGnpBUyrJxEvVgI+1;
	end
	always@(posedge rd_clk or negedge rst)
	begin
		if(!rst)
			nQAnZVgoKyprBQAdRCfA<=0;
		else if(rst_syn)
			nQAnZVgoKyprBQAdRCfA<=0;
		else if(wEtGDzRjafclnvKxgCSP&&nQAnZVgoKyprBQAdRCfA)  
			nQAnZVgoKyprBQAdRCfA<=0;
		else if(one_codeblock_over)
			nQAnZVgoKyprBQAdRCfA<=1;
	end
	always@(posedge rd_clk or negedge rst)
	begin
		if(!rst)
			wEtGDzRjafclnvKxgCSP<=0;
		else if(gStNdqadtalDMswfRuqW==PASS_OVER)
			wEtGDzRjafclnvKxgCSP<=1;            
		else if(flush_over||nQAnZVgoKyprBQAdRCfA)
			wEtGDzRjafclnvKxgCSP<=0;
	end

	always@(posedge wr_clk or negedge rst)
	begin
		if(!rst)
			tQSdMsmQOoDjgNvoiCmq<=0;
		else if(rst_syn)
			tQSdMsmQOoDjgNvoiCmq<=0;
		else if(one_codeblock_over)
			tQSdMsmQOoDjgNvoiCmq<=zero_plane_number; 
	    else if(flush_over)
			tQSdMsmQOoDjgNvoiCmq<=zero_plane_number;
	end

	always@(*)
	begin
	    case(XWSDWJpZwWFziLcqAlai)
 			0:LrLbKGgLtBSEzbICsDNb=DnfnMYzlPFszZtXlGDhW;
    		1:LrLbKGgLtBSEzbICsDNb=NhvFLRUduFzxNErEsMee;
    		2:LrLbKGgLtBSEzbICsDNb=FGUJmfBLDaAxYUKmfnyF;
			default:LrLbKGgLtBSEzbICsDNb=0;
		endcase
	end
	always@(posedge wr_clk or negedge rst)
	begin
	    if(!rst)
		begin
			DnfnMYzlPFszZtXlGDhW <=0;
			NhvFLRUduFzxNErEsMee <=0;
			FGUJmfBLDaAxYUKmfnyF <=0;
		end
		else if(rst_syn)
		begin
			DnfnMYzlPFszZtXlGDhW <=0;
			NhvFLRUduFzxNErEsMee <=0;
			FGUJmfBLDaAxYUKmfnyF <=0;
		end

		else if(flush_over)
		begin
			DnfnMYzlPFszZtXlGDhW <=word_last_flag_plane_sp;
			NhvFLRUduFzxNErEsMee <=word_last_flag_plane_mp;
			FGUJmfBLDaAxYUKmfnyF <=word_last_flag_plane_cp;
		end
	end

	
	
	
	
	always@(*)
	begin
	    if(jMCVmjFKEszeMFGJPhDT)
		begin
			case(lram_address_wr)   
				480:qgkpXRmlTwkWNutDGWMM=MNhKBwmQfBNRRoCGsGYL  ;//{{{
				479:qgkpXRmlTwkWNutDGWMM=CZUlnpSgUmTCmXxNawKq  ;
				478:qgkpXRmlTwkWNutDGWMM=GCKDpTZdSkziHIHQTHTY  ;
				477:qgkpXRmlTwkWNutDGWMM=TbggffYtMBhiLSACnOtm  ;
				476:qgkpXRmlTwkWNutDGWMM=QMFreKPqLMtYHbzgqBQA  ;
				475:qgkpXRmlTwkWNutDGWMM=NlcVQzrrHSpHBCrquBjt  ;
				474:qgkpXRmlTwkWNutDGWMM=FSYqURbHbEaesQcTkdrx  ;
				473:qgkpXRmlTwkWNutDGWMM=qEtkygphCMCbDqrWtklY  ;
				472:qgkpXRmlTwkWNutDGWMM=TLjaqwEsoHtrvWTBQRsK  ;
				471:qgkpXRmlTwkWNutDGWMM=cYsREsbuuQNtJwVuIQtc ;
				470:qgkpXRmlTwkWNutDGWMM=IADijSHmLDuBqTQJOxSa ;
				469:qgkpXRmlTwkWNutDGWMM=BhAYLsocIYeStsZZVTUF ;
				468:qgkpXRmlTwkWNutDGWMM=WQWSkTgEaMFMXPEsFHwg ;
				467:qgkpXRmlTwkWNutDGWMM=WVikipTMfwFUtPMyACXK ;
				466:qgkpXRmlTwkWNutDGWMM=dXrKEPxqSBOppMxaytbW ;
				465:qgkpXRmlTwkWNutDGWMM=NnjJwuwNoVWroSgcnSsE ;
				464:qgkpXRmlTwkWNutDGWMM=ASCWICejFoBbZHMJMVyD ;
				463:qgkpXRmlTwkWNutDGWMM=twyoccXqjNTyiiCHZKgQ ;
				462:qgkpXRmlTwkWNutDGWMM=xvRCARkQSEXoZFEiGfjC ;
				461:qgkpXRmlTwkWNutDGWMM=JjLGddxBYbYmoYBVjdju ;
				460:qgkpXRmlTwkWNutDGWMM=xyvvBnpUfpnejSAdOrIU ;
				459:qgkpXRmlTwkWNutDGWMM=LNWqJGCGvJkqDqnyFdST ;
				458:qgkpXRmlTwkWNutDGWMM=XXnujvRmwKtqZZbYXNom ;
				457:qgkpXRmlTwkWNutDGWMM=rdgcYAhdMEGqsgkVVhHB ;
				456:qgkpXRmlTwkWNutDGWMM=bcCzAdPYbGFOdbqFGtNY ;
				455:qgkpXRmlTwkWNutDGWMM=MRTHuncHaQWNXrTdnjLu ;
				454:qgkpXRmlTwkWNutDGWMM=ZqxWPnvGQEisPGNSDkWt ;
				453:qgkpXRmlTwkWNutDGWMM=jLboxjBIZGftrbnYaDHz ;
				452:qgkpXRmlTwkWNutDGWMM=XPHrltKlkTYeddIYErlL ;
				451:qgkpXRmlTwkWNutDGWMM=DwnEuDbYEGceHCFfntWU ;
				450:qgkpXRmlTwkWNutDGWMM=AhXRxsizDLdrPCSJbgvu ;
				449:qgkpXRmlTwkWNutDGWMM=dRLKJNMhCWjmYIXyBBMS ;
				448:qgkpXRmlTwkWNutDGWMM=qKakmPsWXvxWDjopwmhd ;
				447:qgkpXRmlTwkWNutDGWMM=OfKBQrlHgohHRFQMqPuX ;
				446:qgkpXRmlTwkWNutDGWMM=OMUVfbzXJtBmpgGUlWIN ;
				445:qgkpXRmlTwkWNutDGWMM=pRjKNldSGgrOVpMtRdhl ;
				444:qgkpXRmlTwkWNutDGWMM=FzItXojZYuRrQPYroXqa ;
				443:qgkpXRmlTwkWNutDGWMM=tiASKMApdODRGubKCrIk ;
				442:qgkpXRmlTwkWNutDGWMM=AofWIQWGCHGeAWxyBSnX ;
				441:qgkpXRmlTwkWNutDGWMM=BVZJHRZIRDJUNzlhOXNj ;
				440:qgkpXRmlTwkWNutDGWMM=MJngMbRNrQAqZKOoJbfA ;
				439:qgkpXRmlTwkWNutDGWMM=LKEbaiUcnUkcdhTlxIWn ;
				438:qgkpXRmlTwkWNutDGWMM=PIdKWDjIZqdVETXVKUyz ;
				437:qgkpXRmlTwkWNutDGWMM=TeweoifYlvYAXegPEOev ;
				436:qgkpXRmlTwkWNutDGWMM=aHdPRBehEsBXhVSVEVGI ;
				435:qgkpXRmlTwkWNutDGWMM=EHDzFoGEUiKMcpmeZndO ;
				434:qgkpXRmlTwkWNutDGWMM=iGWdFxfLkcoPAfSnTRiW ;
				433:qgkpXRmlTwkWNutDGWMM=OgwvxakMlGIDTjsTTTrF ;
				432:qgkpXRmlTwkWNutDGWMM=hweOwCSFFCFpnLABsNDz ;
				431:qgkpXRmlTwkWNutDGWMM=kFILldZgHWqtwHcEyrEz ;
				430:qgkpXRmlTwkWNutDGWMM=BHxWpRKaPloRmedcGnVS ;
				429:qgkpXRmlTwkWNutDGWMM=jEDhTzjvJVSeQkYxJusx ;
				428:qgkpXRmlTwkWNutDGWMM=nVWwCingLJiAmNkXNBse ;
				427:qgkpXRmlTwkWNutDGWMM=hdQpCNCsCpWxWjyDHYIf ;
				426:qgkpXRmlTwkWNutDGWMM=mYfjBwhqQaPjGDGuVzVT ;
				425:qgkpXRmlTwkWNutDGWMM=sPdTjZhZROmcYPkfxnHK ;
				424:qgkpXRmlTwkWNutDGWMM=VOSkkJBkJQjLTSFCXXZG ;
				423:qgkpXRmlTwkWNutDGWMM=wnDMhVWFcihAknOuJWgt ;
				422:qgkpXRmlTwkWNutDGWMM=ZJYNMlOSJujZtBMVfIcG ;
				421:qgkpXRmlTwkWNutDGWMM=cUQgUjrarAoCxWvadhrh ;
				420:qgkpXRmlTwkWNutDGWMM=ayPBmMeTERtfSkylBBkl ;
				419:qgkpXRmlTwkWNutDGWMM=zjiIArXGbkjgPxxXfPxg ;
				418:qgkpXRmlTwkWNutDGWMM=YERHnxdykgyyioNNZJSQ ;
				417:qgkpXRmlTwkWNutDGWMM=rNuBwbgCniYGlSgOMCnE ;
				416:qgkpXRmlTwkWNutDGWMM=VjtVxkxLZrdVPkMsyEqe ;
				415:qgkpXRmlTwkWNutDGWMM=fFwIafFNLTVTiIeJUZOi ;
				414:qgkpXRmlTwkWNutDGWMM=JofSpHHAILpRCvnGOmzf ;
				413:qgkpXRmlTwkWNutDGWMM=OeYMhMfjeDdvkecHiLUT ;
				412:qgkpXRmlTwkWNutDGWMM=tVOTCptQSOpsjFBXiksw ;
				411:qgkpXRmlTwkWNutDGWMM=AhXuWEaSPuUvIcwDuFWr ;
				410:qgkpXRmlTwkWNutDGWMM=ekQuaIqPJyasZNSLaQOo ;
				409:qgkpXRmlTwkWNutDGWMM=osvtoSWcIuWcmvZruLsS ;
				408:qgkpXRmlTwkWNutDGWMM=BzXYfwLRzqKLxtfxvmZC ;
				407:qgkpXRmlTwkWNutDGWMM=tgVDzxwqtPquEcvdvFrC ;
				406:qgkpXRmlTwkWNutDGWMM=DzNsyDbNrzFrSyvQMHnd ;
				405:qgkpXRmlTwkWNutDGWMM=iOnjZhBOoaDLaXXeVrwx ;
				404:qgkpXRmlTwkWNutDGWMM=XwvNGtBVJXErWQRUuqBI ;
				403:qgkpXRmlTwkWNutDGWMM=JJgTPGsdUTcAdufkeJgK ;
				402:qgkpXRmlTwkWNutDGWMM=TfnRFMUqcGKfwYVkrOcp ;
				401:qgkpXRmlTwkWNutDGWMM=kuHTqKTEGHJGjcgKEkCF ;
				400:qgkpXRmlTwkWNutDGWMM=FfvTBiXNEwWARzrRMUYh ;
				399:qgkpXRmlTwkWNutDGWMM=VMfdRrsDolDymeMDbscN ;
				398:qgkpXRmlTwkWNutDGWMM=iPuXoTiWLBGZVYAHGaYO ;
				397:qgkpXRmlTwkWNutDGWMM=BaxkmTikPlEanrOALJQn ;
				396:qgkpXRmlTwkWNutDGWMM=TGPYgdsEOqsHqlpqyhVp ;
				395:qgkpXRmlTwkWNutDGWMM=VZaWDekOPjcbcuLkmTCK ;
				394:qgkpXRmlTwkWNutDGWMM=ceSSpUnFGIqusvzAQYyv ;
				393:qgkpXRmlTwkWNutDGWMM=KkgZHqKRoBphLNurbXZv ;
				392:qgkpXRmlTwkWNutDGWMM=BVfKHJmimWhfvhFZYdJC ;
				391:qgkpXRmlTwkWNutDGWMM=XWIoNGOmiUqZuWDNerJA ;
				390:qgkpXRmlTwkWNutDGWMM=ymZNoaOSvkuMNFrKCZJc ;
				389:qgkpXRmlTwkWNutDGWMM=JtPboWbpZfxqTBEEDYyf ;
				388:qgkpXRmlTwkWNutDGWMM=NIzOkTmOrsmtdJpYgwkn ;
				387:qgkpXRmlTwkWNutDGWMM=HPBVjcjYzqThfAZsuBko ;
				386:qgkpXRmlTwkWNutDGWMM=RtOUSNvLjifycdHERnsH ;
				385:qgkpXRmlTwkWNutDGWMM=RHqjRVMUmlsTYhhiTxqt ;
				384:qgkpXRmlTwkWNutDGWMM=irQWRPjnSymTgyEWfOeV ;
				383:qgkpXRmlTwkWNutDGWMM=gHMMxJFDpgQtSoSKsfzc ;
				382:qgkpXRmlTwkWNutDGWMM=XrXzzUeQwqtdbHighLXh ;
				381:qgkpXRmlTwkWNutDGWMM=VXesUOJyNaYiksaASUmr;
				380:qgkpXRmlTwkWNutDGWMM=MjDYzSbWZYtgtBPeFxFX;
				379:qgkpXRmlTwkWNutDGWMM=QocIghyhzPXBoGjaFxEW;
				378:qgkpXRmlTwkWNutDGWMM=aNNRDAQndlQbuwTNoeBC;
				377:qgkpXRmlTwkWNutDGWMM=ganwYnOuHsVFGlnGQGGf;
				376:qgkpXRmlTwkWNutDGWMM=TmUIbPULspEIyexiGCHU;
				375:qgkpXRmlTwkWNutDGWMM=GrWFHsoruHLBTofZiNlc;
				374:qgkpXRmlTwkWNutDGWMM=HemnvXRItkGWOQQBARSS;
				373:qgkpXRmlTwkWNutDGWMM=crDvxwhExTyEkehZAJBR;
				372:qgkpXRmlTwkWNutDGWMM=vqFRiEdZYIvaYIjwIZPo;
				371:qgkpXRmlTwkWNutDGWMM=RiyBtzLqNImqdjYXxYLF;
				370:qgkpXRmlTwkWNutDGWMM=QAZelRxmduKrKymXyprg;
				369:qgkpXRmlTwkWNutDGWMM=IixlIEeyecDFQCcIcXFK;
				368:qgkpXRmlTwkWNutDGWMM=CahtEzYLkeeOsdRKBvoI;
				367:qgkpXRmlTwkWNutDGWMM=hXvwCaJPKLmTlGnIqShO;
				366:qgkpXRmlTwkWNutDGWMM=ZapMeflJnJGQFrDdnzZx;
				365:qgkpXRmlTwkWNutDGWMM=tEZVPsZbWePhmBDkYbkW;
				364:qgkpXRmlTwkWNutDGWMM=VKIhSekuVtyFcvuoBpZH;
				363:qgkpXRmlTwkWNutDGWMM=HHissIgZPvjjCfGzZWgP;
				362:qgkpXRmlTwkWNutDGWMM=ZthEdVQnyODdQJpzqpDX;
				361:qgkpXRmlTwkWNutDGWMM=ZvVAYFyMKYuJjjuLlssM;
				360:qgkpXRmlTwkWNutDGWMM=BDVfxjBZqdgfpcXaqSxS;
				359:qgkpXRmlTwkWNutDGWMM=SYPrSAmIZhepjzRpfAbW;
				358:qgkpXRmlTwkWNutDGWMM=bheecNbLIfuKFYksBrvM;
				357:qgkpXRmlTwkWNutDGWMM=LoFfmBmHEBmQlYvRihJx;
				356:qgkpXRmlTwkWNutDGWMM=RAqkMVQdcCkZqHQrYhTY;
				355:qgkpXRmlTwkWNutDGWMM=JwazcQrhGdLokRSxMIPy;
				354:qgkpXRmlTwkWNutDGWMM=NHwKTvStgXGxecepjZCb;
				353:qgkpXRmlTwkWNutDGWMM=iFhOAEkrfnWgTHHMCrAr;
				352:qgkpXRmlTwkWNutDGWMM=KoZvZIhKhWDYlgwhYWfH;
				351:qgkpXRmlTwkWNutDGWMM=xqkVQlUmzixmBBOWsogM;
				350:qgkpXRmlTwkWNutDGWMM=mZcXpTwcGpwcsXaAXzJZ;
				349:qgkpXRmlTwkWNutDGWMM=tBkJHywSnDHjCloeCKQN;
				348:qgkpXRmlTwkWNutDGWMM=rtIOwgMybhKPbMtTkPHH;
				347:qgkpXRmlTwkWNutDGWMM=ULvOWCBpLiqodnUiPZne;
				346:qgkpXRmlTwkWNutDGWMM=UeCtXzcgpZHmscgLWNgU;
				345:qgkpXRmlTwkWNutDGWMM=NchYslfTwDoJDaIhKQld;
				344:qgkpXRmlTwkWNutDGWMM=vdLrgmXBDTPmGWwCZgJK;
				343:qgkpXRmlTwkWNutDGWMM=fypmfZbmWDbDCXEismjU;
				342:qgkpXRmlTwkWNutDGWMM=FEgAuSjALENQXZOiGFUZ;
				341:qgkpXRmlTwkWNutDGWMM=hUaTrhFAshrngFoHaXaJ;
				340:qgkpXRmlTwkWNutDGWMM=avmhenqBbGIfSBAIabaF;
				339:qgkpXRmlTwkWNutDGWMM=IlmCWYrxdJVqIQywKmAF;
				338:qgkpXRmlTwkWNutDGWMM=GXKZdRvGRyUFWKyHVAFD;
				337:qgkpXRmlTwkWNutDGWMM=PExEfPxznaZHuROUSmfc;
				336:qgkpXRmlTwkWNutDGWMM=DoWtmJCIdGMmwEInsyhi;
				335:qgkpXRmlTwkWNutDGWMM=AtkWXjDVDEZLaumbWZzI;
				334:qgkpXRmlTwkWNutDGWMM=HvOvrGAvaPTzYsRxiQFa;
				333:qgkpXRmlTwkWNutDGWMM=rwPuhbqaLGfEsTZJaDhF;
				332:qgkpXRmlTwkWNutDGWMM=YphfuswJNWiAbvgWEfjm;
				331:qgkpXRmlTwkWNutDGWMM=YhTJCIYfjiXccwQDAncB;
				330:qgkpXRmlTwkWNutDGWMM=KaDxyGuuayhqIxIwbGQG;
				329:qgkpXRmlTwkWNutDGWMM=SCcERabQMmiRZhSuKFqS;
				328:qgkpXRmlTwkWNutDGWMM=ASVDnraQDtLQhInOEyVK;
				327:qgkpXRmlTwkWNutDGWMM=RzDedJWchbeEickgtFOM;
				326:qgkpXRmlTwkWNutDGWMM=qBWQIFhDbnPbANWZJPUR;
				325:qgkpXRmlTwkWNutDGWMM=ONSywhEkLUpjhsBVzOEr;
				324:qgkpXRmlTwkWNutDGWMM=SiWXyZwStCTfnlFxLPQx;
				323:qgkpXRmlTwkWNutDGWMM=ljlzMOdncFtIKCHtOsVQ;
				322:qgkpXRmlTwkWNutDGWMM=sBtkXBZAHFHDVqMZHZdd;
				321:qgkpXRmlTwkWNutDGWMM=ZNywgghYzvszBznGurzE;
				320:qgkpXRmlTwkWNutDGWMM=giByCXZhzRJrKpUfJiYx;
				319:qgkpXRmlTwkWNutDGWMM=NOzoIRcSVgyFREyzzHqs;
				318:qgkpXRmlTwkWNutDGWMM=hvcttLppSPcVixtVRHqN;
				317:qgkpXRmlTwkWNutDGWMM=NXURaWZymtMESRzASoml;
				316:qgkpXRmlTwkWNutDGWMM=OGJwXjhBDuVzMrVxGthI;
				315:qgkpXRmlTwkWNutDGWMM=tDHSWWPwhDHPIdkjEtEW;
				314:qgkpXRmlTwkWNutDGWMM=spPgPLHCbVgdzOmJFakw;
				313:qgkpXRmlTwkWNutDGWMM=NCLfdSDEGhGvIWQaIuMS;
				312:qgkpXRmlTwkWNutDGWMM=NfdfbTCtNjYFDeLLecMe;
				311:qgkpXRmlTwkWNutDGWMM=xIHGyzqgFJSHmjAJEkTk;
				310:qgkpXRmlTwkWNutDGWMM=ffdnbvLvbNGfaiXRKcYD;
				309:qgkpXRmlTwkWNutDGWMM=dDkKlvBKHVNSwGZicnzg;
				308:qgkpXRmlTwkWNutDGWMM=sTYRbAXFBXVNlExKcFRO;
				307:qgkpXRmlTwkWNutDGWMM=QYcegkQFzbKFzvlPxGeR;
				306:qgkpXRmlTwkWNutDGWMM=WCbGOTtDaZUdMPlupDBN;
				305:qgkpXRmlTwkWNutDGWMM=kNoeoxFOMGDTBbVzHlLM;
				304:qgkpXRmlTwkWNutDGWMM=pcsafTpJQiyaKivHSiiO;
				303:qgkpXRmlTwkWNutDGWMM=HhgKJaIdyWwhlApPzTKC;
				302:qgkpXRmlTwkWNutDGWMM=LgxgHDHmFYbeGgXVWgvC;
				301:qgkpXRmlTwkWNutDGWMM=cKBOWdNoOXhznBHdAwlu;
				300:qgkpXRmlTwkWNutDGWMM=KASZraJCWhbAUtfwnLfk;
				299:qgkpXRmlTwkWNutDGWMM=AGPbOkqoDAYNiAUBxYWb;
				298:qgkpXRmlTwkWNutDGWMM=QePGiiHhRVKoAUkzEcSD;
				297:qgkpXRmlTwkWNutDGWMM=ULkqQHcjawmJPPtzcPCS;
				296:qgkpXRmlTwkWNutDGWMM=gVMkJmsMEYFtEfiuwaKj;
				295:qgkpXRmlTwkWNutDGWMM=yHFGaozymIVZZMqtzLDd;
				294:qgkpXRmlTwkWNutDGWMM=XyhfMHNDiNoQgejMGALx;
				293:qgkpXRmlTwkWNutDGWMM=zWhpxSLccsmBmQBUhbQT;
				292:qgkpXRmlTwkWNutDGWMM=xKWgakKpWyTQyBrwYCIS;
				291:qgkpXRmlTwkWNutDGWMM=UkOdSdYxtcxumOakhLgx;
				290:qgkpXRmlTwkWNutDGWMM=nhnBLnxptnOVgbmRStCU;
				289:qgkpXRmlTwkWNutDGWMM=UmXpnIjWZNlfEPEYcDTn;
				288:qgkpXRmlTwkWNutDGWMM=deblhPqNAplcidEXSGqw;
				287:qgkpXRmlTwkWNutDGWMM=GgkZJHLDkhyFsCCzuqLa;
				286:qgkpXRmlTwkWNutDGWMM=pKDUrDrLLWTOdoUxvsyF;
				285:qgkpXRmlTwkWNutDGWMM=JrQYFpYwpBTANpnTvLiU;
				284:qgkpXRmlTwkWNutDGWMM=KencLjTnnSFqjwbVxqJg;
				283:qgkpXRmlTwkWNutDGWMM=TXuaPuUIuhCkLiMhEKiF;
				282:qgkpXRmlTwkWNutDGWMM=aAhmLslHTfVKwKSRWVtp;
				281:qgkpXRmlTwkWNutDGWMM=NJEYMnPHSmEVDftsqzQE;
				280:qgkpXRmlTwkWNutDGWMM=ByBgtRovBsKUVHUQEzwk;
				279:qgkpXRmlTwkWNutDGWMM=pcCSuYOgcgRTEfyKANVf;
				278:qgkpXRmlTwkWNutDGWMM=OOJGXLeAUSSWDwWKvqMN;
				277:qgkpXRmlTwkWNutDGWMM=xzObOtBnVrtyMpWImLGp;
				276:qgkpXRmlTwkWNutDGWMM=fPvbFzCudNRdKXFIwPTW;
				275:qgkpXRmlTwkWNutDGWMM=UCBlEpPTGRkqheRhrmew;
				274:qgkpXRmlTwkWNutDGWMM=rxGiYeZlkdsRNUfrmDKO;
				273:qgkpXRmlTwkWNutDGWMM=BRDRPJjxjaVvUmeEcabW;
				272:qgkpXRmlTwkWNutDGWMM=twevQhSVcRXlOWMZGHZH;
				271:qgkpXRmlTwkWNutDGWMM=hsPTsFDtcTjmyeddHGwC;
				270:qgkpXRmlTwkWNutDGWMM=SnXYHdlnJsKNjOCDlAdk;
				269:qgkpXRmlTwkWNutDGWMM=fzPjNCWXNlBXDEixcMfx;
				268:qgkpXRmlTwkWNutDGWMM=MzxTqhCibhKKovZUinvJ;
				267:qgkpXRmlTwkWNutDGWMM=UjBCIuRFDGUvCwBBwjtv;
				266:qgkpXRmlTwkWNutDGWMM=WLvkMHkFFjSeXeCMFLqU;
				265:qgkpXRmlTwkWNutDGWMM=OdXRCGgZgKmtknFfVeGS;
				264:qgkpXRmlTwkWNutDGWMM=YTagschVaYsVmCoZyGxw;
				263:qgkpXRmlTwkWNutDGWMM=uBDeqwBeWjkFnJPifZac;
				262:qgkpXRmlTwkWNutDGWMM=ChqdVbAPIMvlcdCLZFDM;
				261:qgkpXRmlTwkWNutDGWMM=xVhIWQmsjbKYhycXOZZj;
				260:qgkpXRmlTwkWNutDGWMM=moXSbLoysxSoGKFutzbo;
				259:qgkpXRmlTwkWNutDGWMM=pFrrbOJSlADGwICgxTdA;
				258:qgkpXRmlTwkWNutDGWMM=eFKOOLSSWbJGsojVvoDI;
				257:qgkpXRmlTwkWNutDGWMM=CjkyDsWsnyjeHKnTfjoz;
				256:qgkpXRmlTwkWNutDGWMM=ikgPtqNHSxOonFiPgvOK;
				255:qgkpXRmlTwkWNutDGWMM=JzYgxPBzYqfsNCHdKwWT;
				254:qgkpXRmlTwkWNutDGWMM=rYlFPAhuURCPKCloqLOG;
				253:qgkpXRmlTwkWNutDGWMM=PQEjeJZSeiJdTNkqSiiS;
				252:qgkpXRmlTwkWNutDGWMM=MSaMrnCOKHvvWjrvrLVh;
				251:qgkpXRmlTwkWNutDGWMM=bZovfeygdcHHRKfkxfHl;
				250:qgkpXRmlTwkWNutDGWMM=ATkQsyvByLEkPXEmCGoF;
				249:qgkpXRmlTwkWNutDGWMM=uBtJXFukNYPqTHWppmdv;
				248:qgkpXRmlTwkWNutDGWMM=soNzOmONAzHkpLFWdCtg;
				247:qgkpXRmlTwkWNutDGWMM=lLJeyDbtTaFvkSfqLcWK;
				246:qgkpXRmlTwkWNutDGWMM=lMFLPXTVXadwnVsRrAPI;
				245:qgkpXRmlTwkWNutDGWMM=WPsXEglrQBPoHLKokyap;
				244:qgkpXRmlTwkWNutDGWMM=RqjRxpMaojbkWLGINNMj;
				243:qgkpXRmlTwkWNutDGWMM=CcpgUvVvfmeEoXXGYlgz;
				242:qgkpXRmlTwkWNutDGWMM=yNeJpDTKbQScFfOFsIMP;
				241:qgkpXRmlTwkWNutDGWMM=uVWYpFOIjqHtdFWqJLJL;
				240:qgkpXRmlTwkWNutDGWMM=vCLJZIRyvOOZpamupbmS;
				239:qgkpXRmlTwkWNutDGWMM=JiRCGeWXVDSjvohYatoO;
				238:qgkpXRmlTwkWNutDGWMM=JXVeYnVHSdAGpxmDHgjf;
				237:qgkpXRmlTwkWNutDGWMM=iXlLoGyimBUgUkjZoGvT;
				236:qgkpXRmlTwkWNutDGWMM=JrBVZVJGLbQlQIuxVRMO;
				235:qgkpXRmlTwkWNutDGWMM=MZLrRshlRErhPsqJeccP;
				234:qgkpXRmlTwkWNutDGWMM=KddqRkJXVvlRHkpsKNQL;
				233:qgkpXRmlTwkWNutDGWMM=eKWoIeUrKiPbRIhuWEla;
				232:qgkpXRmlTwkWNutDGWMM=JRsyUSbxyBGBNdlJquOD;
				231:qgkpXRmlTwkWNutDGWMM=mobFFnIZQLEDGamGRCMQ;
				230:qgkpXRmlTwkWNutDGWMM=MIfRQTaujrTsVSIdukaO;
				229:qgkpXRmlTwkWNutDGWMM=qQxKziPkMaoHyxLiZQNv;
				228:qgkpXRmlTwkWNutDGWMM=SbGofGNBnFvEqTbzCMDT;
				227:qgkpXRmlTwkWNutDGWMM=eAyuUdQDmhsyVqUkrWtf;
				226:qgkpXRmlTwkWNutDGWMM=xcrfMbSpXdXRmlkuZRPx;
				225:qgkpXRmlTwkWNutDGWMM=BKSeIpcsVISDrrWyloru;
				224:qgkpXRmlTwkWNutDGWMM=cFxrUFXVhwbgFamPfIXu;
				223:qgkpXRmlTwkWNutDGWMM=EawSFufNSOZZHKtrbfDb;
				222:qgkpXRmlTwkWNutDGWMM=TtHHtKtzZHIcJuWziTSX;
				221:qgkpXRmlTwkWNutDGWMM=KAQFclKTjvNuQpWZONVn;
				220:qgkpXRmlTwkWNutDGWMM=zdDIxzPkCVYUHKycUMxS;
				219:qgkpXRmlTwkWNutDGWMM=yRWhBghWQtDlHOXzOKHV;
				218:qgkpXRmlTwkWNutDGWMM=xzEZrlRsvTQMlJcdcoBA;
				217:qgkpXRmlTwkWNutDGWMM=omKttYZtWwSNmJfXmNhw;
				216:qgkpXRmlTwkWNutDGWMM=TJsrTmKBrLuIryymjrla;
				215:qgkpXRmlTwkWNutDGWMM=UQIvtuLZLyNrLBcITiBh;
				214:qgkpXRmlTwkWNutDGWMM=dewJijMNQrULKORvfOPu;
				213:qgkpXRmlTwkWNutDGWMM=fFCHqQnaXGJtQcWhDHoo;
				212:qgkpXRmlTwkWNutDGWMM=lDVujeiDOsfmAcgTJEeH;
				211:qgkpXRmlTwkWNutDGWMM=tHYVLHNrDsWBBiksZJSh;
				210:qgkpXRmlTwkWNutDGWMM=YGcrryHhhucPWCRpoXpV;
				209:qgkpXRmlTwkWNutDGWMM=vhaFurczuHuVJndQizpm;
				208:qgkpXRmlTwkWNutDGWMM=bAUZnBUzAeFxTBCaAwBD;
				207:qgkpXRmlTwkWNutDGWMM=SJSSeEtWLefcHjjHknTt;
				206:qgkpXRmlTwkWNutDGWMM=RrXElmqzMleQDmHbRetu;
				205:qgkpXRmlTwkWNutDGWMM=RiwCfvabTaSgTyqQQkNP;
				204:qgkpXRmlTwkWNutDGWMM=ijLmWvKcGWYkfmVliDIH;
				203:qgkpXRmlTwkWNutDGWMM=JhZCVmRnYDVfDuTgaJBq;
				202:qgkpXRmlTwkWNutDGWMM=MmtedWLnvMwKkqgwBoYk;
				201:qgkpXRmlTwkWNutDGWMM=xNONPhZsuWCOqfHyKvVw;
				200:qgkpXRmlTwkWNutDGWMM=UYtsWPGzDLbsLPHFFzpM;
				199:qgkpXRmlTwkWNutDGWMM=HaIozTBrCuKZJRqUpAty;
				198:qgkpXRmlTwkWNutDGWMM=ihhBdoTzqImqsCjVxwKM;
				197:qgkpXRmlTwkWNutDGWMM=LPKCNZYNtyFJTUiKvFKI;
				196:qgkpXRmlTwkWNutDGWMM=VcDzTcOFndjUjhnRfxTN;
				195:qgkpXRmlTwkWNutDGWMM=ScSvdbbLcbwcpTKFudIt;
				194:qgkpXRmlTwkWNutDGWMM=ZFOGopcNcymIuYXsiiRw;
				193:qgkpXRmlTwkWNutDGWMM=zVAojGgdEwSIpPjTZZId;
				192:qgkpXRmlTwkWNutDGWMM=qwGWpRzKYsDLRvxcxAAH;
				191:qgkpXRmlTwkWNutDGWMM=WPkpODdzyINGGhuwZyoF;
				190:qgkpXRmlTwkWNutDGWMM=BaxiLnGgFxSKHVKkEWrL;
				189:qgkpXRmlTwkWNutDGWMM=cChsgcLGnvNEmegZREam;
				188:qgkpXRmlTwkWNutDGWMM=FRCWHcmIuMUUWgdYMzWu;
				187:qgkpXRmlTwkWNutDGWMM=QDYrIGBlnoXdNCUflHOP;
				186:qgkpXRmlTwkWNutDGWMM=zzYTnLgksIjwqZSweXMf;
				185:qgkpXRmlTwkWNutDGWMM=cWljGAlocPwsnrDyMjHO;
				184:qgkpXRmlTwkWNutDGWMM=JPYOnWGSGjFuHZfQBaEZ;
				183:qgkpXRmlTwkWNutDGWMM=VzfYJEwelHYPMpUSDmsC;
				182:qgkpXRmlTwkWNutDGWMM=XYQGKDohhXYVCeaCtmre;
				181:qgkpXRmlTwkWNutDGWMM=GbajCDnxXLGTStnsYsds;
				180:qgkpXRmlTwkWNutDGWMM=THlQvXwjkuLqdcMtPxBy;
				179:qgkpXRmlTwkWNutDGWMM=avkJIgYNFpvoyRkxaMTC;
				178:qgkpXRmlTwkWNutDGWMM=yhgnNUWIhVDlrtUDGEZn;
				177:qgkpXRmlTwkWNutDGWMM=lHvULbFfwhQgtqfjhwzH;
				176:qgkpXRmlTwkWNutDGWMM=TymwlUFeZUaLhFoWTZzU;
				175:qgkpXRmlTwkWNutDGWMM=obAWtmAwdFBYPXQlSuSy;
				174:qgkpXRmlTwkWNutDGWMM=VBJGcheVZYcxGpvcuBoi;
				173:qgkpXRmlTwkWNutDGWMM=NpcOSbiIpOcdgCjboENs;
				172:qgkpXRmlTwkWNutDGWMM=PiHYPPmDrZQNPnlqBFSt;
				171:qgkpXRmlTwkWNutDGWMM=rOXoAhCRFHntxISYSkye;
				170:qgkpXRmlTwkWNutDGWMM=IsXHeZVJKogNnFFfJwvx;
				169:qgkpXRmlTwkWNutDGWMM=BtfuDWbiQheMoNKySKtm;
				168:qgkpXRmlTwkWNutDGWMM=lsMUeaCgYLjCPUiUXaIc;
				167:qgkpXRmlTwkWNutDGWMM=kTdnGvNmLrhbepFdhZCh;
				166:qgkpXRmlTwkWNutDGWMM=vKbnovNlLRioZoJsQunL;
				165:qgkpXRmlTwkWNutDGWMM=nXBrtwwgIArkXUbHKAye;
				164:qgkpXRmlTwkWNutDGWMM=czvIYhYPaYPpRHUBJMFc;
				163:qgkpXRmlTwkWNutDGWMM=nsezjQWxmqwzmxCwosDv;
				162:qgkpXRmlTwkWNutDGWMM=ruIyZIesSthmxIaXEtrJ;
				161:qgkpXRmlTwkWNutDGWMM=cXQjLxPFTWRBhlJmdxUJ;
				160:qgkpXRmlTwkWNutDGWMM=GPoMmfciZsakCXuJMdbD;
				159:qgkpXRmlTwkWNutDGWMM=sZUCFycPxeatsZozmHJN;
				158:qgkpXRmlTwkWNutDGWMM=XbnmwpButuNSkogDlbQb;
				157:qgkpXRmlTwkWNutDGWMM=wdkDXnIkWnpQMmswGQeU;
				156:qgkpXRmlTwkWNutDGWMM=KpEHEcApUpQBvCLoAeYT;
				155:qgkpXRmlTwkWNutDGWMM=KsaghLmgaRvpRfCktbJZ;
				154:qgkpXRmlTwkWNutDGWMM=lZVGNfUlVmsuLbJxnQDA;
				153:qgkpXRmlTwkWNutDGWMM=rMBkqrLcKhflEMUYxGkE;
				152:qgkpXRmlTwkWNutDGWMM=wMlYFxkSbZTCTvhQOIei;
				151:qgkpXRmlTwkWNutDGWMM=WQGVbnQQZGQWVmpcxvbb;
				150:qgkpXRmlTwkWNutDGWMM=AzsKalhmBYUitbArLbcU;
				149:qgkpXRmlTwkWNutDGWMM=ekrMWzROxYoWtRpdbLZH;
				148:qgkpXRmlTwkWNutDGWMM=uLMmObkZiwzDlReqMwJN;
				147:qgkpXRmlTwkWNutDGWMM=eAEEsZkRTlfXOeEdICRO;
				146:qgkpXRmlTwkWNutDGWMM=DyXCiZssIzbywKGAbIwY;
				145:qgkpXRmlTwkWNutDGWMM=wBOVUPcFUWzhOUKDlJVa;
				144:qgkpXRmlTwkWNutDGWMM=BCsgCSHvysHWLteqbRMX;
				143:qgkpXRmlTwkWNutDGWMM=FrvVghZEElOfAJGPEURk;
				142:qgkpXRmlTwkWNutDGWMM=DHNpdfPdlvcIeMhPYCBD;
				141:qgkpXRmlTwkWNutDGWMM=ByKBiFClfZeeoBwNqVdH;
				140:qgkpXRmlTwkWNutDGWMM=muXlkjUrAqYazTUUGcVg;
				139:qgkpXRmlTwkWNutDGWMM=rZlIolWetZZffpSrlMAn;
				138:qgkpXRmlTwkWNutDGWMM=fCxfzzVrwjVhwiuAOpOD;
				137:qgkpXRmlTwkWNutDGWMM=VHDrEEGVFWccsKXzbEjD;
				136:qgkpXRmlTwkWNutDGWMM=pgbmZFwAnGMkExuHZexG;
				135:qgkpXRmlTwkWNutDGWMM=CYTIFZXRYHDOwAOpYhTY;
				134:qgkpXRmlTwkWNutDGWMM=hzujftnKaamrwjRBenpS;
				133:qgkpXRmlTwkWNutDGWMM=DwBiXGPwomcqrFUiwGKO;
				132:qgkpXRmlTwkWNutDGWMM=TxOTbaXnfvTWWAEMVKsT;
				131:qgkpXRmlTwkWNutDGWMM=VBPMSBgUzhZWqifRFXLt;
				130:qgkpXRmlTwkWNutDGWMM=fBEMznDkaUpJbucpUFUs;
				129:qgkpXRmlTwkWNutDGWMM=RXuUWWKfwotmzMaIdOHs;
				128:qgkpXRmlTwkWNutDGWMM=DScSrBltRCaJuMKRHxjp;
				127:qgkpXRmlTwkWNutDGWMM=yKhNJjIQvjuuxuKGtNvD;
				126:qgkpXRmlTwkWNutDGWMM=MBLbhXLxXGZHZERKIoYb;
				125:qgkpXRmlTwkWNutDGWMM=AiFthZhNPfZiXSnyPCOt;
				124:qgkpXRmlTwkWNutDGWMM=uDpYTElkHJsWMgegRIkv;
				123:qgkpXRmlTwkWNutDGWMM=LqJHECWMJlDdyFDTTZZH;
				122:qgkpXRmlTwkWNutDGWMM=ohfsyAOCKLVNdUfnlZGT;
				121:qgkpXRmlTwkWNutDGWMM=MOoDdDePAGBzQbLCZlwX;
				120:qgkpXRmlTwkWNutDGWMM=MHLazVdHgoSmGTltAxsJ;
				119:qgkpXRmlTwkWNutDGWMM=CYSqcBzpHDXSSATrgQjL;
				118:qgkpXRmlTwkWNutDGWMM=rPKZMoWgFDpDSJXXQmEU;
				117:qgkpXRmlTwkWNutDGWMM=hniufLGfdzmHbDIvsTIo;
				116:qgkpXRmlTwkWNutDGWMM=wTfPVycgpDcgGCOQhJjH;
				115:qgkpXRmlTwkWNutDGWMM=lcOMvsbHZmIJccXoDkqZ;
				114:qgkpXRmlTwkWNutDGWMM=UKirjTCurmcGUGGogrnh;
				113:qgkpXRmlTwkWNutDGWMM=KVLRCNcgwgdezgxdbtiz;
				112:qgkpXRmlTwkWNutDGWMM=ISUkQBFCDDhkmXDnEdVT;
				111:qgkpXRmlTwkWNutDGWMM=wLiUXxuAUdxCuAoAbUxH;
				110:qgkpXRmlTwkWNutDGWMM=vQNMUmgdbJJDFKzsjqLK;
				109:qgkpXRmlTwkWNutDGWMM=PPaVHoPQXNFqYDIgCroQ;
				108:qgkpXRmlTwkWNutDGWMM=fZmgOJpwMcdeRjEcecxZ;
				107:qgkpXRmlTwkWNutDGWMM=pXxRQDEgUJLwgwAsNvmV;
				106:qgkpXRmlTwkWNutDGWMM=JWyFVCrskBwarfgMzbIK;
				105:qgkpXRmlTwkWNutDGWMM=nLMIykvKsueQiebJRjaB;
				104:qgkpXRmlTwkWNutDGWMM=MwUAnLVNdEpwKFXarSrE;
				103:qgkpXRmlTwkWNutDGWMM=rwKFeNNlWzDutFvKudZd;
				102:qgkpXRmlTwkWNutDGWMM=YFTuhpacOohGrtlEUgyn;
				101:qgkpXRmlTwkWNutDGWMM=orsjfJIPQQvjIhvrnfZT;
				100:qgkpXRmlTwkWNutDGWMM=beooHOrejCcWcSXDuAMs;
				99 :qgkpXRmlTwkWNutDGWMM=wLFqLqnhtGKyjhXVaXLu;
				98 :qgkpXRmlTwkWNutDGWMM=VhlEwlgxfirfMpIAJZhE;
				97 :qgkpXRmlTwkWNutDGWMM=ybSCwixJTEhXYyRpEeDj;
				96 :qgkpXRmlTwkWNutDGWMM=PLAwknGzfcioZVaFOQCX;
				95 :qgkpXRmlTwkWNutDGWMM=WdDdHRBJZdBPCxmYbWdk;
				94 :qgkpXRmlTwkWNutDGWMM=BIxIzsQvWljjGYxMCQtS;
				93 :qgkpXRmlTwkWNutDGWMM=TZYUrtPvAdyOAezlYVJO;
				92 :qgkpXRmlTwkWNutDGWMM=qPqZhRZBobhmAXNGrsmh;
				91 :qgkpXRmlTwkWNutDGWMM=BCGaGkllXBcyohBosHqS;
				90 :qgkpXRmlTwkWNutDGWMM=pcgiabuotmBHXKOYDDAq;
				89 :qgkpXRmlTwkWNutDGWMM=VidvAsXIfsppEpKtZeYc;
				88 :qgkpXRmlTwkWNutDGWMM=lGfaCxQtDihDBzWEuyaH;
				87 :qgkpXRmlTwkWNutDGWMM=ucwrtDfHQDZIjkmTmCvN;
				86 :qgkpXRmlTwkWNutDGWMM=dayIzRpYaQRnEjXynbCm;
				85 :qgkpXRmlTwkWNutDGWMM=vqgpItmCwuhiwKZyFXMt;
				84 :qgkpXRmlTwkWNutDGWMM=FnVEwsGKlXZfUqxZGqHn;
				83 :qgkpXRmlTwkWNutDGWMM=bitnzrgsExKEWSXnsRZq;
				82 :qgkpXRmlTwkWNutDGWMM=eYsNwIgUOqnSppAZBKfW;
				81 :qgkpXRmlTwkWNutDGWMM=FXTNpbkOJRifihZRkFUk;
				80 :qgkpXRmlTwkWNutDGWMM=UCyPKegIVHgIqztViRHP;
				79 :qgkpXRmlTwkWNutDGWMM=urwbynurHojveDuzQAqY;
				78 :qgkpXRmlTwkWNutDGWMM=djsdiJHbeUEoOocTIVAL;
				77 :qgkpXRmlTwkWNutDGWMM=juEeWiBDxjlSPOBoDWca;
				76 :qgkpXRmlTwkWNutDGWMM=ZfhQiwfaJoKgwqVVBKhf;
				75 :qgkpXRmlTwkWNutDGWMM=SNnVNrhdPUfxhixiespl;
				74 :qgkpXRmlTwkWNutDGWMM=cHHoYqPSIzoxFEuXvNLY;
				73 :qgkpXRmlTwkWNutDGWMM=hLpCUWbILJOjqbDhVEwn;
				72 :qgkpXRmlTwkWNutDGWMM=itXQCyFacJzvPyzfGwVe;
				71 :qgkpXRmlTwkWNutDGWMM=iujmIQQClXPYAKjueUBD;
				70 :qgkpXRmlTwkWNutDGWMM=BjdcbpGuKPxnpZzFTfte;
				69 :qgkpXRmlTwkWNutDGWMM=ZQFzyLJsVraTCGkqQcZA;
				68 :qgkpXRmlTwkWNutDGWMM=fADZyEOwTyWvSQFgOnwG;
				67 :qgkpXRmlTwkWNutDGWMM=xbhqvpXrDTlnyBNQeAlC;
				66 :qgkpXRmlTwkWNutDGWMM=usigvHtlPqTHmByMEGLy;
				65 :qgkpXRmlTwkWNutDGWMM=EqRnSoIxQaLPlCNmpBmq;
				64 :qgkpXRmlTwkWNutDGWMM=VzsEzvUFwafgXDXiMnOI;
				63 :qgkpXRmlTwkWNutDGWMM=qjQChEpAPSbKmoDGRppN;
				62 :qgkpXRmlTwkWNutDGWMM=XBdmfGxuWrXGMBFOANKF;
				61 :qgkpXRmlTwkWNutDGWMM=iHWmgCopJntOccGPObxn;
				60 :qgkpXRmlTwkWNutDGWMM=eeoTbTyuwxPCsjuUGnLj;
				59 :qgkpXRmlTwkWNutDGWMM=MkxrURKJtUzHVTfBwhoO;
				58 :qgkpXRmlTwkWNutDGWMM=USFkaPtDBVOjbGpLXKUX;
				57 :qgkpXRmlTwkWNutDGWMM=xcBSpPXNgyeMCKwBcsxX;
				56 :qgkpXRmlTwkWNutDGWMM=APZhwjfiYOuKluWEaTIj;
				55 :qgkpXRmlTwkWNutDGWMM=eiYeGwmYgODBCzcNuNtn;
				54 :qgkpXRmlTwkWNutDGWMM=rmoQVcRSrSeskIibJzCc;
				53 :qgkpXRmlTwkWNutDGWMM=AzSDmFqniQGEkrUvtcQd;
				52 :qgkpXRmlTwkWNutDGWMM=BYQMYRDRDKXGHnLYQyKL;
				51 :qgkpXRmlTwkWNutDGWMM=iYaojeeenaSObFkfIEyS;
				50 :qgkpXRmlTwkWNutDGWMM=OvjWCALXGQonpSVNSUDx;
				49 :qgkpXRmlTwkWNutDGWMM=QNSQONiKmlvpucXZsAKo;
				48 :qgkpXRmlTwkWNutDGWMM=RKLbOFQSgMkwEdftvnBQ;
				47 :qgkpXRmlTwkWNutDGWMM=hoPvrLDkwXFTkYESCUcp;
				46 :qgkpXRmlTwkWNutDGWMM=hShwACbdYktXmGxyazAM;
				45 :qgkpXRmlTwkWNutDGWMM=puehHutFkvCRvoGqbSYp;
				44 :qgkpXRmlTwkWNutDGWMM=CSpvXCVkXjBnWvAFEiDG;
				43 :qgkpXRmlTwkWNutDGWMM=GBnbMGmdJLNqPHpTRJqo;
				42 :qgkpXRmlTwkWNutDGWMM=PQFlqUWXvhfFTKRniEDA;
				41 :qgkpXRmlTwkWNutDGWMM=mNQfwTdWpUOnxIhbTYfU;
				40 :qgkpXRmlTwkWNutDGWMM=ldQowZgtPeXlzjFcyWQl;
				39 :qgkpXRmlTwkWNutDGWMM=HYWHYpKWyjTHzWIzGNeE;
				38 :qgkpXRmlTwkWNutDGWMM=vsHmuANStIQsYgoNHsHw;
				37 :qgkpXRmlTwkWNutDGWMM=tYWmIUymjXADFjUmKFpP;
				36 :qgkpXRmlTwkWNutDGWMM=OQmggBTvOqhAXBiDJeaP;
				35 :qgkpXRmlTwkWNutDGWMM=EFcUAERFHbivPwgHAMQa;
				34 :qgkpXRmlTwkWNutDGWMM=jpbydIYGKyCwhjgemImi;
				33 :qgkpXRmlTwkWNutDGWMM=OVYjPuZDVHOTTeuFPkrT;
				32 :qgkpXRmlTwkWNutDGWMM=DqhwOfIUxBzsVSgEjWzC;
				31 :qgkpXRmlTwkWNutDGWMM=plztNCDwyKBliboMvXKs;
				30 :qgkpXRmlTwkWNutDGWMM=GojVETmCGfWcYwVYimBv;
				29 :qgkpXRmlTwkWNutDGWMM=aogDiFiAXQqphSrsQbJV;
				28 :qgkpXRmlTwkWNutDGWMM=rCOKgSoVLfXaUWFdsBnJ;
				27 :qgkpXRmlTwkWNutDGWMM=ZuONZDcmHxALaUULMEAA;
				26 :qgkpXRmlTwkWNutDGWMM=KIjEeYrBOSrzUMqGYBsV;
				25 :qgkpXRmlTwkWNutDGWMM=ZBocacKljeyYorCiQgzQ;
				24 :qgkpXRmlTwkWNutDGWMM=mqazMnBgYnlLqLRzaNYx;
				23 :qgkpXRmlTwkWNutDGWMM=oyfKvpCwkpoCCxTglCJr;
				22 :qgkpXRmlTwkWNutDGWMM=NGNEGckWnRLaqnjOKOmx;
				21 :qgkpXRmlTwkWNutDGWMM=cVWqyzzrUUodYFbrorBz;
				20 :qgkpXRmlTwkWNutDGWMM=RjwugczIYXEQzzmUrnYh;
				19 :qgkpXRmlTwkWNutDGWMM=lEqWgKBWIbLvYwrXeDtN;
				18 :qgkpXRmlTwkWNutDGWMM=DhnZhzYLzUMXzuxLMdpR;
				17 :qgkpXRmlTwkWNutDGWMM=WwogGcAbNuwPRaXHfllR;
				16 :qgkpXRmlTwkWNutDGWMM=fymbKnqnRYaHIRuPXxle;
				15 :qgkpXRmlTwkWNutDGWMM=nJWkhXEkUmrasSyMThpL;
				14 :qgkpXRmlTwkWNutDGWMM=qXNWBYTrrKKKGSroThrT;
				13 :qgkpXRmlTwkWNutDGWMM=OWgmvdYcTEmvwkEuDkJS;
				12 :qgkpXRmlTwkWNutDGWMM=urpaOisfjSiDXEZoTBsG;
				11 :qgkpXRmlTwkWNutDGWMM=mveotDylkopgLZJFFBVl;
				10 :qgkpXRmlTwkWNutDGWMM=CCXECvtOeIBEOFePtIRw;
				9  :qgkpXRmlTwkWNutDGWMM=iYYwLjjGMjLikfxxrxIB;
				8  :qgkpXRmlTwkWNutDGWMM=BJhcDugYXUoZuTXYBzJg;
				7  :qgkpXRmlTwkWNutDGWMM=wpEZHrezpouBVvAiIOpn;
				6  :qgkpXRmlTwkWNutDGWMM=omjfRcaEwaSdXWjgQYUv;
				5  :qgkpXRmlTwkWNutDGWMM=aWXCrpICnOAsyXgkDTDT;
				4  :qgkpXRmlTwkWNutDGWMM=HjXRkNnhDmrrYeoZLfga;
				3  :qgkpXRmlTwkWNutDGWMM=zDWiKpAenkhcNZIBSNiT;
				2  :qgkpXRmlTwkWNutDGWMM=UfyNbuBOwMXEdumKnlqN;
				1  :qgkpXRmlTwkWNutDGWMM=LYSwVHbgNGVrAkuDLmxY;
				0  :qgkpXRmlTwkWNutDGWMM=0;//}}}
				default:qgkpXRmlTwkWNutDGWMM=0;
			endcase
		end
		else qgkpXRmlTwkWNutDGWMM=0;
	end
	
	always@(posedge rd_clk or negedge rst)
	begin
	    if(!rst)
			GVfnzKKftzXfxeBqPQMD<=0;
		else if(rst_syn)
			GVfnzKKftzXfxeBqPQMD<=0;
		else if(jMCVmjFKEszeMFGJPhDT)  
		begin
			GVfnzKKftzXfxeBqPQMD<=GVfnzKKftzXfxeBqPQMD+qgkpXRmlTwkWNutDGWMM;
		end
	end
	
	
	always@(*)
	begin
	    case(compression_ratio)
			0:target_byte_number=4919 ;
			1:target_byte_number=2458  ;
			2:target_byte_number=1229  ;
			3:target_byte_number=614   ;
			4:target_byte_number=307   ;
			default:target_byte_number=0;
	    endcase
	end
	always@(posedge rd_clk or negedge rst)
	begin
	    if(!rst)
			lram_write_en<=0;
		else if(rst_syn)
			lram_write_en<=0;
		else if((gStNdqadtalDMswfRuqW==SHIFT_PASS_SECOND_HEADER)||(gStNdqadtalDMswfRuqW==SHIFT_CODESTREAM)||(gStNdqadtalDMswfRuqW==SHIFT_PASS_FIRST_HEADER)||(gStNdqadtalDMswfRuqW==SHIFT_OVER_FLAG))
			lram_write_en<=1;
		else lram_write_en<=0;
	end
	
	always@(posedge wr_clk)
	begin
	    XmWQfEltjOUqcNLDCtfd<=one_codeblock_over;
		pyhAjCtAJLKGgXMclzgY<=XmWQfEltjOUqcNLDCtfd;
		MPFTDVkljwqlROSuxXcP<=pyhAjCtAJLKGgXMclzgY;
	end
	
	always@(*)
	begin
		if(eojmGbYrZBcDvhuhplcn)
		begin
			case(XWSDWJpZwWFziLcqAlai)
				0:aSItvOfWsSQOkHOHMzuM=iGrqtIPPBFPUhGunhSdw;
    			1:aSItvOfWsSQOkHOHMzuM=CZceBwenUmhgWecdrVuw;
    			2:aSItvOfWsSQOkHOHMzuM=FODhltaveISdQIJPBJhJ;
				default:aSItvOfWsSQOkHOHMzuM=0;
			endcase
		end
		else
		begin
			case(XWSDWJpZwWFziLcqAlai)
				0:aSItvOfWsSQOkHOHMzuM=mBUfUweOiYOTkxaNfvqZ;
    			1:aSItvOfWsSQOkHOHMzuM=XCEBnusbPkduEdkiHxFK;
    			2:aSItvOfWsSQOkHOHMzuM=UKLUuuVquDsMMMMhkoJV;
				default:aSItvOfWsSQOkHOHMzuM=0;
			endcase
		end
	end
	
	always@(*)
	begin
	    case(gStNdqadtalDMswfRuqW)
			 CAL_SLOPE_1:ESEFEoPuTgYdvrsaqlOz=rczbRGCFDOHKNTiwObwc[37:8];
			 CAL_SLOPE_2:ESEFEoPuTgYdvrsaqlOz=OHenhlDjGfxNrcoKTDTe[37:8];
			 default:ESEFEoPuTgYdvrsaqlOz=0;
			endcase
	end
	
	always@(*)
	begin
	    casex(ESEFEoPuTgYdvrsaqlOz)
			30'b1x_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=29;
			30'b01_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=28;
			30'b00_1xxx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=27;
			30'b00_01xx_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=26;
			30'b00_001x_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=25;
			30'b00_0001_xxxx_xxxx_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=24;
			30'b00_0000_1xxx_xxxx_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=23;
			30'b00_0000_01xx_xxxx_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=22;
			30'b00_0000_001x_xxxx_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=21;
			30'b00_0000_0001_xxxx_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=20;
			30'b00_0000_0000_1xxx_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=19;
			30'b00_0000_0000_01xx_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=18;
			30'b00_0000_0000_001x_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=17;
			30'b00_0000_0000_0001_xxxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=16;
			30'b00_0000_0000_0000_1xxx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=15;
			30'b00_0000_0000_0000_01xx_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=14;
			30'b00_0000_0000_0000_001x_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=13;
			30'b00_0000_0000_0000_0001_xxxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=12;
			30'b00_0000_0000_0000_0000_1xxx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=11;
			30'b00_0000_0000_0000_0000_01xx_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT=10;
			30'b00_0000_0000_0000_0000_001x_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT= 9;
			30'b00_0000_0000_0000_0000_0001_xxxx_xxxx:ARQLJGuTZBnFJHXDoAkT= 8;
			30'b00_0000_0000_0000_0000_0000_1xxx_xxxx:ARQLJGuTZBnFJHXDoAkT= 7;
			30'b00_0000_0000_0000_0000_0000_01xx_xxxx:ARQLJGuTZBnFJHXDoAkT= 6;
			30'b00_0000_0000_0000_0000_0000_001x_xxxx:ARQLJGuTZBnFJHXDoAkT= 5;
			30'b00_0000_0000_0000_0000_0000_0001_xxxx:ARQLJGuTZBnFJHXDoAkT= 4;
			30'b00_0000_0000_0000_0000_0000_0000_1xxx:ARQLJGuTZBnFJHXDoAkT= 3;
			30'b00_0000_0000_0000_0000_0000_0000_01xx:ARQLJGuTZBnFJHXDoAkT= 2;
			30'b00_0000_0000_0000_0000_0000_0000_001x:ARQLJGuTZBnFJHXDoAkT= 1;
			30'b00_0000_0000_0000_0000_0000_0000_0001:ARQLJGuTZBnFJHXDoAkT= 0;
			30'b00_0000_0000_0000_0000_0000_0000_0000:ARQLJGuTZBnFJHXDoAkT= 0;
			default:ARQLJGuTZBnFJHXDoAkT= 5'bx;
			endcase
		
	end

	
	always@(posedge rd_clk or negedge rst)
	begin
	    if(!rst)
		begin
			MNhKBwmQfBNRRoCGsGYL  <=0;//{{{
			CZUlnpSgUmTCmXxNawKq  <=0;
			GCKDpTZdSkziHIHQTHTY  <=0;
			TbggffYtMBhiLSACnOtm  <=0;
			QMFreKPqLMtYHbzgqBQA  <=0;
			NlcVQzrrHSpHBCrquBjt  <=0;
			FSYqURbHbEaesQcTkdrx  <=0;
			qEtkygphCMCbDqrWtklY  <=0;
			TLjaqwEsoHtrvWTBQRsK  <=0;
			cYsREsbuuQNtJwVuIQtc <=0;
			IADijSHmLDuBqTQJOxSa <=0;
			BhAYLsocIYeStsZZVTUF <=0;
			WQWSkTgEaMFMXPEsFHwg <=0;
			WVikipTMfwFUtPMyACXK <=0;
			dXrKEPxqSBOppMxaytbW <=0;
			NnjJwuwNoVWroSgcnSsE <=0;
			ASCWICejFoBbZHMJMVyD <=0;
			twyoccXqjNTyiiCHZKgQ <=0;
			xvRCARkQSEXoZFEiGfjC <=0;
			JjLGddxBYbYmoYBVjdju <=0;
			xyvvBnpUfpnejSAdOrIU <=0;
			LNWqJGCGvJkqDqnyFdST <=0;
			XXnujvRmwKtqZZbYXNom <=0;
			rdgcYAhdMEGqsgkVVhHB <=0;
			bcCzAdPYbGFOdbqFGtNY <=0;
			MRTHuncHaQWNXrTdnjLu <=0;
			ZqxWPnvGQEisPGNSDkWt <=0;
			jLboxjBIZGftrbnYaDHz <=0;
			XPHrltKlkTYeddIYErlL <=0;
			DwnEuDbYEGceHCFfntWU <=0;
			AhXRxsizDLdrPCSJbgvu <=0;
			dRLKJNMhCWjmYIXyBBMS <=0;
			qKakmPsWXvxWDjopwmhd <=0;
			OfKBQrlHgohHRFQMqPuX <=0;
			OMUVfbzXJtBmpgGUlWIN <=0;
			pRjKNldSGgrOVpMtRdhl <=0;
			FzItXojZYuRrQPYroXqa <=0;
			tiASKMApdODRGubKCrIk <=0;
			AofWIQWGCHGeAWxyBSnX <=0;
			BVZJHRZIRDJUNzlhOXNj <=0;
			MJngMbRNrQAqZKOoJbfA <=0;
			LKEbaiUcnUkcdhTlxIWn <=0;
			PIdKWDjIZqdVETXVKUyz <=0;
			TeweoifYlvYAXegPEOev <=0;
			aHdPRBehEsBXhVSVEVGI <=0;
			EHDzFoGEUiKMcpmeZndO <=0;
			iGWdFxfLkcoPAfSnTRiW <=0;
			OgwvxakMlGIDTjsTTTrF <=0;
			hweOwCSFFCFpnLABsNDz <=0;
			kFILldZgHWqtwHcEyrEz <=0;
			BHxWpRKaPloRmedcGnVS <=0;
			jEDhTzjvJVSeQkYxJusx <=0;
			nVWwCingLJiAmNkXNBse <=0;
			hdQpCNCsCpWxWjyDHYIf <=0;
			mYfjBwhqQaPjGDGuVzVT <=0;
			sPdTjZhZROmcYPkfxnHK <=0;
			VOSkkJBkJQjLTSFCXXZG <=0;
			wnDMhVWFcihAknOuJWgt <=0;
			ZJYNMlOSJujZtBMVfIcG <=0;
			cUQgUjrarAoCxWvadhrh <=0;
			ayPBmMeTERtfSkylBBkl <=0;
			zjiIArXGbkjgPxxXfPxg <=0;
			YERHnxdykgyyioNNZJSQ <=0;
			rNuBwbgCniYGlSgOMCnE <=0;
			VjtVxkxLZrdVPkMsyEqe <=0;
			fFwIafFNLTVTiIeJUZOi <=0;
			JofSpHHAILpRCvnGOmzf <=0;
			OeYMhMfjeDdvkecHiLUT <=0;
			tVOTCptQSOpsjFBXiksw <=0;
			AhXuWEaSPuUvIcwDuFWr <=0;
			ekQuaIqPJyasZNSLaQOo <=0;
			osvtoSWcIuWcmvZruLsS <=0;
			BzXYfwLRzqKLxtfxvmZC <=0;
			tgVDzxwqtPquEcvdvFrC <=0;
			DzNsyDbNrzFrSyvQMHnd <=0;
			iOnjZhBOoaDLaXXeVrwx <=0;
			XwvNGtBVJXErWQRUuqBI <=0;
			JJgTPGsdUTcAdufkeJgK <=0;
			TfnRFMUqcGKfwYVkrOcp <=0;
			kuHTqKTEGHJGjcgKEkCF <=0;
			FfvTBiXNEwWARzrRMUYh <=0;
			VMfdRrsDolDymeMDbscN <=0;
			iPuXoTiWLBGZVYAHGaYO <=0;
			BaxkmTikPlEanrOALJQn <=0;
			TGPYgdsEOqsHqlpqyhVp <=0;
			VZaWDekOPjcbcuLkmTCK <=0;
			ceSSpUnFGIqusvzAQYyv <=0;
			KkgZHqKRoBphLNurbXZv <=0;
			BVfKHJmimWhfvhFZYdJC <=0;
			XWIoNGOmiUqZuWDNerJA <=0;
			ymZNoaOSvkuMNFrKCZJc <=0;
			JtPboWbpZfxqTBEEDYyf <=0;
			NIzOkTmOrsmtdJpYgwkn <=0;
			HPBVjcjYzqThfAZsuBko <=0;
			RtOUSNvLjifycdHERnsH <=0;
			RHqjRVMUmlsTYhhiTxqt <=0;
			irQWRPjnSymTgyEWfOeV <=0;
			gHMMxJFDpgQtSoSKsfzc <=0;
			XrXzzUeQwqtdbHighLXh <=0;
			VXesUOJyNaYiksaASUmr<=0; 
			MjDYzSbWZYtgtBPeFxFX<=0; 
			QocIghyhzPXBoGjaFxEW<=0; 
			aNNRDAQndlQbuwTNoeBC<=0; 
			ganwYnOuHsVFGlnGQGGf<=0; 
			TmUIbPULspEIyexiGCHU<=0; 
			GrWFHsoruHLBTofZiNlc<=0; 
			HemnvXRItkGWOQQBARSS<=0; 
			crDvxwhExTyEkehZAJBR<=0; 
			vqFRiEdZYIvaYIjwIZPo<=0; 
			RiyBtzLqNImqdjYXxYLF<=0; 
			QAZelRxmduKrKymXyprg<=0; 
			IixlIEeyecDFQCcIcXFK<=0; 
			CahtEzYLkeeOsdRKBvoI<=0; 
			hXvwCaJPKLmTlGnIqShO<=0; 
			ZapMeflJnJGQFrDdnzZx<=0; 
			tEZVPsZbWePhmBDkYbkW<=0; 
			VKIhSekuVtyFcvuoBpZH<=0; 
			HHissIgZPvjjCfGzZWgP<=0; 
			ZthEdVQnyODdQJpzqpDX<=0; 
			ZvVAYFyMKYuJjjuLlssM<=0; 
			BDVfxjBZqdgfpcXaqSxS<=0; 
			SYPrSAmIZhepjzRpfAbW<=0; 
			bheecNbLIfuKFYksBrvM<=0; 
			LoFfmBmHEBmQlYvRihJx<=0; 
			RAqkMVQdcCkZqHQrYhTY<=0; 
			JwazcQrhGdLokRSxMIPy<=0; 
			NHwKTvStgXGxecepjZCb<=0; 
			iFhOAEkrfnWgTHHMCrAr<=0; 
			KoZvZIhKhWDYlgwhYWfH<=0; 
			xqkVQlUmzixmBBOWsogM<=0; 
			mZcXpTwcGpwcsXaAXzJZ<=0; 
			tBkJHywSnDHjCloeCKQN<=0; 
			rtIOwgMybhKPbMtTkPHH<=0; 
			ULvOWCBpLiqodnUiPZne<=0; 
			UeCtXzcgpZHmscgLWNgU<=0; 
			NchYslfTwDoJDaIhKQld<=0; 
			vdLrgmXBDTPmGWwCZgJK<=0; 
			fypmfZbmWDbDCXEismjU<=0; 
			FEgAuSjALENQXZOiGFUZ<=0; 
			hUaTrhFAshrngFoHaXaJ<=0; 
			avmhenqBbGIfSBAIabaF<=0; 
			IlmCWYrxdJVqIQywKmAF<=0; 
			GXKZdRvGRyUFWKyHVAFD<=0; 
			PExEfPxznaZHuROUSmfc<=0; 
			DoWtmJCIdGMmwEInsyhi<=0; 
			AtkWXjDVDEZLaumbWZzI<=0; 
			HvOvrGAvaPTzYsRxiQFa<=0; 
			rwPuhbqaLGfEsTZJaDhF<=0; 
			YphfuswJNWiAbvgWEfjm<=0; 
			YhTJCIYfjiXccwQDAncB<=0; 
			KaDxyGuuayhqIxIwbGQG<=0; 
			SCcERabQMmiRZhSuKFqS<=0; 
			ASVDnraQDtLQhInOEyVK<=0; 
			RzDedJWchbeEickgtFOM<=0; 
			qBWQIFhDbnPbANWZJPUR<=0; 
			ONSywhEkLUpjhsBVzOEr<=0; 
			SiWXyZwStCTfnlFxLPQx<=0; 
			ljlzMOdncFtIKCHtOsVQ<=0; 
			sBtkXBZAHFHDVqMZHZdd<=0; 
			ZNywgghYzvszBznGurzE<=0; 
			giByCXZhzRJrKpUfJiYx<=0; 
			NOzoIRcSVgyFREyzzHqs<=0; 
			hvcttLppSPcVixtVRHqN<=0; 
			NXURaWZymtMESRzASoml<=0; 
			OGJwXjhBDuVzMrVxGthI<=0; 
			tDHSWWPwhDHPIdkjEtEW<=0; 
			spPgPLHCbVgdzOmJFakw<=0; 
			NCLfdSDEGhGvIWQaIuMS<=0; 
			NfdfbTCtNjYFDeLLecMe<=0; 
			xIHGyzqgFJSHmjAJEkTk<=0; 
			ffdnbvLvbNGfaiXRKcYD<=0; 
			dDkKlvBKHVNSwGZicnzg<=0; 
			sTYRbAXFBXVNlExKcFRO<=0; 
			QYcegkQFzbKFzvlPxGeR<=0; 
			WCbGOTtDaZUdMPlupDBN<=0; 
			kNoeoxFOMGDTBbVzHlLM<=0; 
			pcsafTpJQiyaKivHSiiO<=0; 
			HhgKJaIdyWwhlApPzTKC<=0; 
			LgxgHDHmFYbeGgXVWgvC<=0; 
			cKBOWdNoOXhznBHdAwlu<=0; 
			KASZraJCWhbAUtfwnLfk<=0; 
			AGPbOkqoDAYNiAUBxYWb<=0; 
			QePGiiHhRVKoAUkzEcSD<=0; 
			ULkqQHcjawmJPPtzcPCS<=0; 
			gVMkJmsMEYFtEfiuwaKj<=0; 
			yHFGaozymIVZZMqtzLDd<=0; 
			XyhfMHNDiNoQgejMGALx<=0; 
			zWhpxSLccsmBmQBUhbQT<=0; 
			xKWgakKpWyTQyBrwYCIS<=0; 
			UkOdSdYxtcxumOakhLgx<=0; 
			nhnBLnxptnOVgbmRStCU<=0; 
			UmXpnIjWZNlfEPEYcDTn<=0; 
			deblhPqNAplcidEXSGqw<=0; 
			GgkZJHLDkhyFsCCzuqLa<=0; 
			pKDUrDrLLWTOdoUxvsyF<=0; 
			JrQYFpYwpBTANpnTvLiU<=0; 
			KencLjTnnSFqjwbVxqJg<=0; 
			TXuaPuUIuhCkLiMhEKiF<=0; 
			aAhmLslHTfVKwKSRWVtp<=0; 
			NJEYMnPHSmEVDftsqzQE<=0; 
			ByBgtRovBsKUVHUQEzwk<=0; 
			pcCSuYOgcgRTEfyKANVf<=0; 
			OOJGXLeAUSSWDwWKvqMN<=0; 
			xzObOtBnVrtyMpWImLGp<=0; 
			fPvbFzCudNRdKXFIwPTW<=0; 
			UCBlEpPTGRkqheRhrmew<=0; 
			rxGiYeZlkdsRNUfrmDKO<=0; 
			BRDRPJjxjaVvUmeEcabW<=0; 
			twevQhSVcRXlOWMZGHZH<=0; 
			hsPTsFDtcTjmyeddHGwC<=0; 
			SnXYHdlnJsKNjOCDlAdk<=0; 
			fzPjNCWXNlBXDEixcMfx<=0; 
			MzxTqhCibhKKovZUinvJ<=0; 
			UjBCIuRFDGUvCwBBwjtv<=0; 
			WLvkMHkFFjSeXeCMFLqU<=0; 
			OdXRCGgZgKmtknFfVeGS<=0; 
			YTagschVaYsVmCoZyGxw<=0; 
			uBDeqwBeWjkFnJPifZac<=0; 
			ChqdVbAPIMvlcdCLZFDM<=0; 
			xVhIWQmsjbKYhycXOZZj<=0; 
			moXSbLoysxSoGKFutzbo<=0; 
			pFrrbOJSlADGwICgxTdA<=0; 
			eFKOOLSSWbJGsojVvoDI<=0; 
			CjkyDsWsnyjeHKnTfjoz<=0; 
			ikgPtqNHSxOonFiPgvOK<=0; 
			JzYgxPBzYqfsNCHdKwWT<=0; 
			rYlFPAhuURCPKCloqLOG<=0; 
			PQEjeJZSeiJdTNkqSiiS<=0; 
			MSaMrnCOKHvvWjrvrLVh<=0; 
			bZovfeygdcHHRKfkxfHl<=0; 
			ATkQsyvByLEkPXEmCGoF<=0; 
			uBtJXFukNYPqTHWppmdv<=0; 
			soNzOmONAzHkpLFWdCtg<=0; 
			lLJeyDbtTaFvkSfqLcWK<=0; 
			lMFLPXTVXadwnVsRrAPI<=0; 
			WPsXEglrQBPoHLKokyap<=0; 
			RqjRxpMaojbkWLGINNMj<=0; 
			CcpgUvVvfmeEoXXGYlgz<=0; 
			yNeJpDTKbQScFfOFsIMP<=0; 
			uVWYpFOIjqHtdFWqJLJL<=0; 
			vCLJZIRyvOOZpamupbmS<=0; 
			JiRCGeWXVDSjvohYatoO<=0; 
			JXVeYnVHSdAGpxmDHgjf<=0; 
			iXlLoGyimBUgUkjZoGvT<=0; 
			JrBVZVJGLbQlQIuxVRMO<=0; 
			MZLrRshlRErhPsqJeccP<=0; 
			KddqRkJXVvlRHkpsKNQL<=0; 
			eKWoIeUrKiPbRIhuWEla<=0; 
			JRsyUSbxyBGBNdlJquOD<=0; 
			mobFFnIZQLEDGamGRCMQ<=0; 
			MIfRQTaujrTsVSIdukaO<=0; 
			qQxKziPkMaoHyxLiZQNv<=0; 
			SbGofGNBnFvEqTbzCMDT<=0; 
			eAyuUdQDmhsyVqUkrWtf<=0; 
			xcrfMbSpXdXRmlkuZRPx<=0; 
			BKSeIpcsVISDrrWyloru<=0; 
			cFxrUFXVhwbgFamPfIXu<=0; 
			EawSFufNSOZZHKtrbfDb<=0; 
			TtHHtKtzZHIcJuWziTSX<=0; 
			KAQFclKTjvNuQpWZONVn<=0; 
			zdDIxzPkCVYUHKycUMxS<=0; 
			yRWhBghWQtDlHOXzOKHV<=0; 
			xzEZrlRsvTQMlJcdcoBA<=0; 
			omKttYZtWwSNmJfXmNhw<=0; 
			TJsrTmKBrLuIryymjrla<=0; 
			UQIvtuLZLyNrLBcITiBh<=0; 
			dewJijMNQrULKORvfOPu<=0; 
			fFCHqQnaXGJtQcWhDHoo<=0; 
			lDVujeiDOsfmAcgTJEeH<=0; 
			tHYVLHNrDsWBBiksZJSh<=0; 
			YGcrryHhhucPWCRpoXpV<=0; 
			vhaFurczuHuVJndQizpm<=0; 
			bAUZnBUzAeFxTBCaAwBD<=0; 
			SJSSeEtWLefcHjjHknTt<=0; 
			RrXElmqzMleQDmHbRetu<=0; 
			RiwCfvabTaSgTyqQQkNP<=0; 
			ijLmWvKcGWYkfmVliDIH<=0; 
			JhZCVmRnYDVfDuTgaJBq<=0; 
			MmtedWLnvMwKkqgwBoYk<=0; 
			xNONPhZsuWCOqfHyKvVw<=0; 
			UYtsWPGzDLbsLPHFFzpM<=0; 
			HaIozTBrCuKZJRqUpAty<=0; 
			ihhBdoTzqImqsCjVxwKM<=0; 
			LPKCNZYNtyFJTUiKvFKI<=0; 
			VcDzTcOFndjUjhnRfxTN<=0; 
			ScSvdbbLcbwcpTKFudIt<=0; 
			ZFOGopcNcymIuYXsiiRw<=0; 
			zVAojGgdEwSIpPjTZZId<=0; 
			qwGWpRzKYsDLRvxcxAAH<=0; 
			WPkpODdzyINGGhuwZyoF<=0; 
			BaxiLnGgFxSKHVKkEWrL<=0; 
			cChsgcLGnvNEmegZREam<=0; 
			FRCWHcmIuMUUWgdYMzWu<=0; 
			QDYrIGBlnoXdNCUflHOP<=0; 
			zzYTnLgksIjwqZSweXMf<=0; 
			cWljGAlocPwsnrDyMjHO<=0; 
			JPYOnWGSGjFuHZfQBaEZ<=0; 
			VzfYJEwelHYPMpUSDmsC<=0; 
			XYQGKDohhXYVCeaCtmre<=0; 
			GbajCDnxXLGTStnsYsds<=0; 
			THlQvXwjkuLqdcMtPxBy<=0; 
			avkJIgYNFpvoyRkxaMTC<=0; 
			yhgnNUWIhVDlrtUDGEZn<=0; 
			lHvULbFfwhQgtqfjhwzH<=0; 
			TymwlUFeZUaLhFoWTZzU<=0; 
			obAWtmAwdFBYPXQlSuSy<=0; 
			VBJGcheVZYcxGpvcuBoi<=0; 
			NpcOSbiIpOcdgCjboENs<=0; 
			PiHYPPmDrZQNPnlqBFSt<=0; 
			rOXoAhCRFHntxISYSkye<=0; 
			IsXHeZVJKogNnFFfJwvx<=0; 
			BtfuDWbiQheMoNKySKtm<=0; 
			lsMUeaCgYLjCPUiUXaIc<=0; 
			kTdnGvNmLrhbepFdhZCh<=0; 
			vKbnovNlLRioZoJsQunL<=0; 
			nXBrtwwgIArkXUbHKAye<=0; 
			czvIYhYPaYPpRHUBJMFc<=0; 
			nsezjQWxmqwzmxCwosDv<=0; 
			ruIyZIesSthmxIaXEtrJ<=0; 
			cXQjLxPFTWRBhlJmdxUJ<=0; 
			GPoMmfciZsakCXuJMdbD<=0; 
			sZUCFycPxeatsZozmHJN<=0; 
			XbnmwpButuNSkogDlbQb<=0; 
			wdkDXnIkWnpQMmswGQeU<=0; 
			KpEHEcApUpQBvCLoAeYT<=0; 
			KsaghLmgaRvpRfCktbJZ<=0; 
			lZVGNfUlVmsuLbJxnQDA<=0; 
			rMBkqrLcKhflEMUYxGkE<=0; 
			wMlYFxkSbZTCTvhQOIei<=0; 
			WQGVbnQQZGQWVmpcxvbb<=0; 
			AzsKalhmBYUitbArLbcU<=0; 
			ekrMWzROxYoWtRpdbLZH<=0; 
			uLMmObkZiwzDlReqMwJN<=0; 
			eAEEsZkRTlfXOeEdICRO<=0; 
			DyXCiZssIzbywKGAbIwY<=0; 
			wBOVUPcFUWzhOUKDlJVa<=0; 
			BCsgCSHvysHWLteqbRMX<=0; 
			FrvVghZEElOfAJGPEURk<=0; 
			DHNpdfPdlvcIeMhPYCBD<=0; 
			ByKBiFClfZeeoBwNqVdH<=0; 
			muXlkjUrAqYazTUUGcVg<=0; 
			rZlIolWetZZffpSrlMAn<=0; 
			fCxfzzVrwjVhwiuAOpOD<=0; 
			VHDrEEGVFWccsKXzbEjD<=0; 
			pgbmZFwAnGMkExuHZexG<=0; 
			CYTIFZXRYHDOwAOpYhTY<=0; 
			hzujftnKaamrwjRBenpS<=0; 
			DwBiXGPwomcqrFUiwGKO<=0; 
			TxOTbaXnfvTWWAEMVKsT<=0; 
			VBPMSBgUzhZWqifRFXLt<=0; 
			fBEMznDkaUpJbucpUFUs<=0; 
			RXuUWWKfwotmzMaIdOHs<=0; 
			DScSrBltRCaJuMKRHxjp<=0; 
			yKhNJjIQvjuuxuKGtNvD<=0; 
			MBLbhXLxXGZHZERKIoYb<=0; 
			AiFthZhNPfZiXSnyPCOt<=0; 
			uDpYTElkHJsWMgegRIkv<=0; 
			LqJHECWMJlDdyFDTTZZH<=0; 
			ohfsyAOCKLVNdUfnlZGT<=0; 
			MOoDdDePAGBzQbLCZlwX<=0; 
			MHLazVdHgoSmGTltAxsJ<=0; 
			CYSqcBzpHDXSSATrgQjL<=0; 
			rPKZMoWgFDpDSJXXQmEU<=0; 
			hniufLGfdzmHbDIvsTIo<=0; 
			wTfPVycgpDcgGCOQhJjH<=0; 
			lcOMvsbHZmIJccXoDkqZ<=0; 
			UKirjTCurmcGUGGogrnh<=0; 
			KVLRCNcgwgdezgxdbtiz<=0; 
			ISUkQBFCDDhkmXDnEdVT<=0; 
			wLiUXxuAUdxCuAoAbUxH<=0; 
			vQNMUmgdbJJDFKzsjqLK<=0; 
			PPaVHoPQXNFqYDIgCroQ<=0; 
			fZmgOJpwMcdeRjEcecxZ<=0; 
			pXxRQDEgUJLwgwAsNvmV<=0; 
			JWyFVCrskBwarfgMzbIK<=0; 
			nLMIykvKsueQiebJRjaB<=0; 
			MwUAnLVNdEpwKFXarSrE<=0; 
			rwKFeNNlWzDutFvKudZd<=0; 
			YFTuhpacOohGrtlEUgyn<=0; 
			orsjfJIPQQvjIhvrnfZT<=0; 
			beooHOrejCcWcSXDuAMs<=0; 
			wLFqLqnhtGKyjhXVaXLu<=0; 
			VhlEwlgxfirfMpIAJZhE<=0; 
			ybSCwixJTEhXYyRpEeDj<=0; 
			PLAwknGzfcioZVaFOQCX<=0; 
			WdDdHRBJZdBPCxmYbWdk<=0; 
			BIxIzsQvWljjGYxMCQtS<=0; 
			TZYUrtPvAdyOAezlYVJO<=0; 
			qPqZhRZBobhmAXNGrsmh<=0; 
			BCGaGkllXBcyohBosHqS<=0; 
			pcgiabuotmBHXKOYDDAq<=0; 
			VidvAsXIfsppEpKtZeYc<=0; 
			lGfaCxQtDihDBzWEuyaH<=0; 
			ucwrtDfHQDZIjkmTmCvN<=0; 
			dayIzRpYaQRnEjXynbCm<=0; 
			vqgpItmCwuhiwKZyFXMt<=0; 
			FnVEwsGKlXZfUqxZGqHn<=0; 
			bitnzrgsExKEWSXnsRZq<=0; 
			eYsNwIgUOqnSppAZBKfW<=0; 
			FXTNpbkOJRifihZRkFUk<=0; 
			UCyPKegIVHgIqztViRHP<=0; 
			urwbynurHojveDuzQAqY<=0; 
			djsdiJHbeUEoOocTIVAL<=0; 
			juEeWiBDxjlSPOBoDWca<=0; 
			ZfhQiwfaJoKgwqVVBKhf<=0; 
			SNnVNrhdPUfxhixiespl<=0; 
			cHHoYqPSIzoxFEuXvNLY<=0; 
			hLpCUWbILJOjqbDhVEwn<=0; 
			itXQCyFacJzvPyzfGwVe<=0; 
			iujmIQQClXPYAKjueUBD<=0; 
			BjdcbpGuKPxnpZzFTfte<=0; 
			ZQFzyLJsVraTCGkqQcZA<=0; 
			fADZyEOwTyWvSQFgOnwG<=0; 
			xbhqvpXrDTlnyBNQeAlC<=0; 
			usigvHtlPqTHmByMEGLy<=0; 
			EqRnSoIxQaLPlCNmpBmq<=0; 
			VzsEzvUFwafgXDXiMnOI<=0; 
			qjQChEpAPSbKmoDGRppN<=0; 
			XBdmfGxuWrXGMBFOANKF<=0; 
			iHWmgCopJntOccGPObxn<=0; 
			eeoTbTyuwxPCsjuUGnLj<=0; 
			MkxrURKJtUzHVTfBwhoO<=0; 
			USFkaPtDBVOjbGpLXKUX<=0; 
			xcBSpPXNgyeMCKwBcsxX<=0; 
			APZhwjfiYOuKluWEaTIj<=0; 
			eiYeGwmYgODBCzcNuNtn<=0; 
			rmoQVcRSrSeskIibJzCc<=0; 
			AzSDmFqniQGEkrUvtcQd<=0; 
			BYQMYRDRDKXGHnLYQyKL<=0; 
			iYaojeeenaSObFkfIEyS<=0; 
			OvjWCALXGQonpSVNSUDx<=0; 
			QNSQONiKmlvpucXZsAKo<=0; 
			RKLbOFQSgMkwEdftvnBQ<=0; 
			hoPvrLDkwXFTkYESCUcp<=0; 
			hShwACbdYktXmGxyazAM<=0; 
			puehHutFkvCRvoGqbSYp<=0; 
			CSpvXCVkXjBnWvAFEiDG<=0; 
			GBnbMGmdJLNqPHpTRJqo<=0; 
			PQFlqUWXvhfFTKRniEDA<=0; 
			mNQfwTdWpUOnxIhbTYfU<=0; 
			ldQowZgtPeXlzjFcyWQl<=0; 
			HYWHYpKWyjTHzWIzGNeE<=0; 
			vsHmuANStIQsYgoNHsHw<=0; 
			tYWmIUymjXADFjUmKFpP<=0; 
			OQmggBTvOqhAXBiDJeaP<=0; 
			EFcUAERFHbivPwgHAMQa<=0; 
			jpbydIYGKyCwhjgemImi<=0; 
			OVYjPuZDVHOTTeuFPkrT<=0; 
			DqhwOfIUxBzsVSgEjWzC<=0; 
			plztNCDwyKBliboMvXKs<=0; 
			GojVETmCGfWcYwVYimBv<=0; 
			aogDiFiAXQqphSrsQbJV<=0; 
			rCOKgSoVLfXaUWFdsBnJ<=0; 
			ZuONZDcmHxALaUULMEAA<=0; 
			KIjEeYrBOSrzUMqGYBsV<=0; 
			ZBocacKljeyYorCiQgzQ<=0; 
			mqazMnBgYnlLqLRzaNYx<=0; 
			oyfKvpCwkpoCCxTglCJr<=0; 
			NGNEGckWnRLaqnjOKOmx<=0; 
			cVWqyzzrUUodYFbrorBz<=0; 
			RjwugczIYXEQzzmUrnYh<=0; 
			lEqWgKBWIbLvYwrXeDtN<=0; 
			DhnZhzYLzUMXzuxLMdpR<=0; 
			WwogGcAbNuwPRaXHfllR<=0; 
			fymbKnqnRYaHIRuPXxle<=0; 
			nJWkhXEkUmrasSyMThpL<=0; 
			qXNWBYTrrKKKGSroThrT<=0; 
			OWgmvdYcTEmvwkEuDkJS<=0; 
			urpaOisfjSiDXEZoTBsG<=0; 
			mveotDylkopgLZJFFBVl<=0; 
			CCXECvtOeIBEOFePtIRw<=0; 
			iYYwLjjGMjLikfxxrxIB<=0; 
			BJhcDugYXUoZuTXYBzJg<=0; 
			wpEZHrezpouBVvAiIOpn<=0; 
			omjfRcaEwaSdXWjgQYUv<=0; 
			aWXCrpICnOAsyXgkDTDT<=0; 
			HjXRkNnhDmrrYeoZLfga<=0; 
			zDWiKpAenkhcNZIBSNiT<=0; 
			UfyNbuBOwMXEdumKnlqN<=0; 
			LYSwVHbgNGVrAkuDLmxY<=0;
		end
		else if(rst_syn)
		begin
			MNhKBwmQfBNRRoCGsGYL  <=0;
			CZUlnpSgUmTCmXxNawKq  <=0;
			GCKDpTZdSkziHIHQTHTY  <=0;
			TbggffYtMBhiLSACnOtm  <=0;
			QMFreKPqLMtYHbzgqBQA  <=0;
			NlcVQzrrHSpHBCrquBjt  <=0;
			FSYqURbHbEaesQcTkdrx  <=0;
			qEtkygphCMCbDqrWtklY  <=0;
			TLjaqwEsoHtrvWTBQRsK  <=0;
			cYsREsbuuQNtJwVuIQtc <=0;
			IADijSHmLDuBqTQJOxSa <=0;
			BhAYLsocIYeStsZZVTUF <=0;
			WQWSkTgEaMFMXPEsFHwg <=0;
			WVikipTMfwFUtPMyACXK <=0;
			dXrKEPxqSBOppMxaytbW <=0;
			NnjJwuwNoVWroSgcnSsE <=0;
			ASCWICejFoBbZHMJMVyD <=0;
			twyoccXqjNTyiiCHZKgQ <=0;
			xvRCARkQSEXoZFEiGfjC <=0;
			JjLGddxBYbYmoYBVjdju <=0;
			xyvvBnpUfpnejSAdOrIU <=0;
			LNWqJGCGvJkqDqnyFdST <=0;
			XXnujvRmwKtqZZbYXNom <=0;
			rdgcYAhdMEGqsgkVVhHB <=0;
			bcCzAdPYbGFOdbqFGtNY <=0;
			MRTHuncHaQWNXrTdnjLu <=0;
			ZqxWPnvGQEisPGNSDkWt <=0;
			jLboxjBIZGftrbnYaDHz <=0;
			XPHrltKlkTYeddIYErlL <=0;
			DwnEuDbYEGceHCFfntWU <=0;
			AhXRxsizDLdrPCSJbgvu <=0;
			dRLKJNMhCWjmYIXyBBMS <=0;
			qKakmPsWXvxWDjopwmhd <=0;
			OfKBQrlHgohHRFQMqPuX <=0;
			OMUVfbzXJtBmpgGUlWIN <=0;
			pRjKNldSGgrOVpMtRdhl <=0;
			FzItXojZYuRrQPYroXqa <=0;
			tiASKMApdODRGubKCrIk <=0;
			AofWIQWGCHGeAWxyBSnX <=0;
			BVZJHRZIRDJUNzlhOXNj <=0;
			MJngMbRNrQAqZKOoJbfA <=0;
			LKEbaiUcnUkcdhTlxIWn <=0;
			PIdKWDjIZqdVETXVKUyz <=0;
			TeweoifYlvYAXegPEOev <=0;
			aHdPRBehEsBXhVSVEVGI <=0;
			EHDzFoGEUiKMcpmeZndO <=0;
			iGWdFxfLkcoPAfSnTRiW <=0;
			OgwvxakMlGIDTjsTTTrF <=0;
			hweOwCSFFCFpnLABsNDz <=0;
			kFILldZgHWqtwHcEyrEz <=0;
			BHxWpRKaPloRmedcGnVS <=0;
			jEDhTzjvJVSeQkYxJusx <=0;
			nVWwCingLJiAmNkXNBse <=0;
			hdQpCNCsCpWxWjyDHYIf <=0;
			mYfjBwhqQaPjGDGuVzVT <=0;
			sPdTjZhZROmcYPkfxnHK <=0;
			VOSkkJBkJQjLTSFCXXZG <=0;
			wnDMhVWFcihAknOuJWgt <=0;
			ZJYNMlOSJujZtBMVfIcG <=0;
			cUQgUjrarAoCxWvadhrh <=0;
			ayPBmMeTERtfSkylBBkl <=0;
			zjiIArXGbkjgPxxXfPxg <=0;
			YERHnxdykgyyioNNZJSQ <=0;
			rNuBwbgCniYGlSgOMCnE <=0;
			VjtVxkxLZrdVPkMsyEqe <=0;
			fFwIafFNLTVTiIeJUZOi <=0;
			JofSpHHAILpRCvnGOmzf <=0;
			OeYMhMfjeDdvkecHiLUT <=0;
			tVOTCptQSOpsjFBXiksw <=0;
			AhXuWEaSPuUvIcwDuFWr <=0;
			ekQuaIqPJyasZNSLaQOo <=0;
			osvtoSWcIuWcmvZruLsS <=0;
			BzXYfwLRzqKLxtfxvmZC <=0;
			tgVDzxwqtPquEcvdvFrC <=0;
			DzNsyDbNrzFrSyvQMHnd <=0;
			iOnjZhBOoaDLaXXeVrwx <=0;
			XwvNGtBVJXErWQRUuqBI <=0;
			JJgTPGsdUTcAdufkeJgK <=0;
			TfnRFMUqcGKfwYVkrOcp <=0;
			kuHTqKTEGHJGjcgKEkCF <=0;
			FfvTBiXNEwWARzrRMUYh <=0;
			VMfdRrsDolDymeMDbscN <=0;
			iPuXoTiWLBGZVYAHGaYO <=0;
			BaxkmTikPlEanrOALJQn <=0;
			TGPYgdsEOqsHqlpqyhVp <=0;
			VZaWDekOPjcbcuLkmTCK <=0;
			ceSSpUnFGIqusvzAQYyv <=0;
			KkgZHqKRoBphLNurbXZv <=0;
			BVfKHJmimWhfvhFZYdJC <=0;
			XWIoNGOmiUqZuWDNerJA <=0;
			ymZNoaOSvkuMNFrKCZJc <=0;
			JtPboWbpZfxqTBEEDYyf <=0;
			NIzOkTmOrsmtdJpYgwkn <=0;
			HPBVjcjYzqThfAZsuBko <=0;
			RtOUSNvLjifycdHERnsH <=0;
			RHqjRVMUmlsTYhhiTxqt <=0;
			irQWRPjnSymTgyEWfOeV <=0;
			gHMMxJFDpgQtSoSKsfzc <=0;
			XrXzzUeQwqtdbHighLXh <=0;
			VXesUOJyNaYiksaASUmr<=0; 
			MjDYzSbWZYtgtBPeFxFX<=0; 
			QocIghyhzPXBoGjaFxEW<=0; 
			aNNRDAQndlQbuwTNoeBC<=0; 
			ganwYnOuHsVFGlnGQGGf<=0; 
			TmUIbPULspEIyexiGCHU<=0; 
			GrWFHsoruHLBTofZiNlc<=0; 
			HemnvXRItkGWOQQBARSS<=0; 
			crDvxwhExTyEkehZAJBR<=0; 
			vqFRiEdZYIvaYIjwIZPo<=0; 
			RiyBtzLqNImqdjYXxYLF<=0; 
			QAZelRxmduKrKymXyprg<=0; 
			IixlIEeyecDFQCcIcXFK<=0; 
			CahtEzYLkeeOsdRKBvoI<=0; 
			hXvwCaJPKLmTlGnIqShO<=0; 
			ZapMeflJnJGQFrDdnzZx<=0; 
			tEZVPsZbWePhmBDkYbkW<=0; 
			VKIhSekuVtyFcvuoBpZH<=0; 
			HHissIgZPvjjCfGzZWgP<=0; 
			ZthEdVQnyODdQJpzqpDX<=0; 
			ZvVAYFyMKYuJjjuLlssM<=0; 
			BDVfxjBZqdgfpcXaqSxS<=0; 
			SYPrSAmIZhepjzRpfAbW<=0; 
			bheecNbLIfuKFYksBrvM<=0; 
			LoFfmBmHEBmQlYvRihJx<=0; 
			RAqkMVQdcCkZqHQrYhTY<=0; 
			JwazcQrhGdLokRSxMIPy<=0; 
			NHwKTvStgXGxecepjZCb<=0; 
			iFhOAEkrfnWgTHHMCrAr<=0; 
			KoZvZIhKhWDYlgwhYWfH<=0; 
			xqkVQlUmzixmBBOWsogM<=0; 
			mZcXpTwcGpwcsXaAXzJZ<=0; 
			tBkJHywSnDHjCloeCKQN<=0; 
			rtIOwgMybhKPbMtTkPHH<=0; 
			ULvOWCBpLiqodnUiPZne<=0; 
			UeCtXzcgpZHmscgLWNgU<=0; 
			NchYslfTwDoJDaIhKQld<=0; 
			vdLrgmXBDTPmGWwCZgJK<=0; 
			fypmfZbmWDbDCXEismjU<=0; 
			FEgAuSjALENQXZOiGFUZ<=0; 
			hUaTrhFAshrngFoHaXaJ<=0; 
			avmhenqBbGIfSBAIabaF<=0; 
			IlmCWYrxdJVqIQywKmAF<=0; 
			GXKZdRvGRyUFWKyHVAFD<=0; 
			PExEfPxznaZHuROUSmfc<=0; 
			DoWtmJCIdGMmwEInsyhi<=0; 
			AtkWXjDVDEZLaumbWZzI<=0; 
			HvOvrGAvaPTzYsRxiQFa<=0; 
			rwPuhbqaLGfEsTZJaDhF<=0; 
			YphfuswJNWiAbvgWEfjm<=0; 
			YhTJCIYfjiXccwQDAncB<=0; 
			KaDxyGuuayhqIxIwbGQG<=0; 
			SCcERabQMmiRZhSuKFqS<=0; 
			ASVDnraQDtLQhInOEyVK<=0; 
			RzDedJWchbeEickgtFOM<=0; 
			qBWQIFhDbnPbANWZJPUR<=0; 
			ONSywhEkLUpjhsBVzOEr<=0; 
			SiWXyZwStCTfnlFxLPQx<=0; 
			ljlzMOdncFtIKCHtOsVQ<=0; 
			sBtkXBZAHFHDVqMZHZdd<=0; 
			ZNywgghYzvszBznGurzE<=0; 
			giByCXZhzRJrKpUfJiYx<=0; 
			NOzoIRcSVgyFREyzzHqs<=0; 
			hvcttLppSPcVixtVRHqN<=0; 
			NXURaWZymtMESRzASoml<=0; 
			OGJwXjhBDuVzMrVxGthI<=0; 
			tDHSWWPwhDHPIdkjEtEW<=0; 
			spPgPLHCbVgdzOmJFakw<=0; 
			NCLfdSDEGhGvIWQaIuMS<=0; 
			NfdfbTCtNjYFDeLLecMe<=0; 
			xIHGyzqgFJSHmjAJEkTk<=0; 
			ffdnbvLvbNGfaiXRKcYD<=0; 
			dDkKlvBKHVNSwGZicnzg<=0; 
			sTYRbAXFBXVNlExKcFRO<=0; 
			QYcegkQFzbKFzvlPxGeR<=0; 
			WCbGOTtDaZUdMPlupDBN<=0; 
			kNoeoxFOMGDTBbVzHlLM<=0; 
			pcsafTpJQiyaKivHSiiO<=0; 
			HhgKJaIdyWwhlApPzTKC<=0; 
			LgxgHDHmFYbeGgXVWgvC<=0; 
			cKBOWdNoOXhznBHdAwlu<=0; 
			KASZraJCWhbAUtfwnLfk<=0; 
			AGPbOkqoDAYNiAUBxYWb<=0; 
			QePGiiHhRVKoAUkzEcSD<=0; 
			ULkqQHcjawmJPPtzcPCS<=0; 
			gVMkJmsMEYFtEfiuwaKj<=0; 
			yHFGaozymIVZZMqtzLDd<=0; 
			XyhfMHNDiNoQgejMGALx<=0; 
			zWhpxSLccsmBmQBUhbQT<=0; 
			xKWgakKpWyTQyBrwYCIS<=0; 
			UkOdSdYxtcxumOakhLgx<=0; 
			nhnBLnxptnOVgbmRStCU<=0; 
			UmXpnIjWZNlfEPEYcDTn<=0; 
			deblhPqNAplcidEXSGqw<=0; 
			GgkZJHLDkhyFsCCzuqLa<=0; 
			pKDUrDrLLWTOdoUxvsyF<=0; 
			JrQYFpYwpBTANpnTvLiU<=0; 
			KencLjTnnSFqjwbVxqJg<=0; 
			TXuaPuUIuhCkLiMhEKiF<=0; 
			aAhmLslHTfVKwKSRWVtp<=0; 
			NJEYMnPHSmEVDftsqzQE<=0; 
			ByBgtRovBsKUVHUQEzwk<=0; 
			pcCSuYOgcgRTEfyKANVf<=0; 
			OOJGXLeAUSSWDwWKvqMN<=0; 
			xzObOtBnVrtyMpWImLGp<=0; 
			fPvbFzCudNRdKXFIwPTW<=0; 
			UCBlEpPTGRkqheRhrmew<=0; 
			rxGiYeZlkdsRNUfrmDKO<=0; 
			BRDRPJjxjaVvUmeEcabW<=0; 
			twevQhSVcRXlOWMZGHZH<=0; 
			hsPTsFDtcTjmyeddHGwC<=0; 
			SnXYHdlnJsKNjOCDlAdk<=0; 
			fzPjNCWXNlBXDEixcMfx<=0; 
			MzxTqhCibhKKovZUinvJ<=0; 
			UjBCIuRFDGUvCwBBwjtv<=0; 
			WLvkMHkFFjSeXeCMFLqU<=0; 
			OdXRCGgZgKmtknFfVeGS<=0; 
			YTagschVaYsVmCoZyGxw<=0; 
			uBDeqwBeWjkFnJPifZac<=0; 
			ChqdVbAPIMvlcdCLZFDM<=0; 
			xVhIWQmsjbKYhycXOZZj<=0; 
			moXSbLoysxSoGKFutzbo<=0; 
			pFrrbOJSlADGwICgxTdA<=0; 
			eFKOOLSSWbJGsojVvoDI<=0; 
			CjkyDsWsnyjeHKnTfjoz<=0; 
			ikgPtqNHSxOonFiPgvOK<=0; 
			JzYgxPBzYqfsNCHdKwWT<=0; 
			rYlFPAhuURCPKCloqLOG<=0; 
			PQEjeJZSeiJdTNkqSiiS<=0; 
			MSaMrnCOKHvvWjrvrLVh<=0; 
			bZovfeygdcHHRKfkxfHl<=0; 
			ATkQsyvByLEkPXEmCGoF<=0; 
			uBtJXFukNYPqTHWppmdv<=0; 
			soNzOmONAzHkpLFWdCtg<=0; 
			lLJeyDbtTaFvkSfqLcWK<=0; 
			lMFLPXTVXadwnVsRrAPI<=0; 
			WPsXEglrQBPoHLKokyap<=0; 
			RqjRxpMaojbkWLGINNMj<=0; 
			CcpgUvVvfmeEoXXGYlgz<=0; 
			yNeJpDTKbQScFfOFsIMP<=0; 
			uVWYpFOIjqHtdFWqJLJL<=0; 
			vCLJZIRyvOOZpamupbmS<=0; 
			JiRCGeWXVDSjvohYatoO<=0; 
			JXVeYnVHSdAGpxmDHgjf<=0; 
			iXlLoGyimBUgUkjZoGvT<=0; 
			JrBVZVJGLbQlQIuxVRMO<=0; 
			MZLrRshlRErhPsqJeccP<=0; 
			KddqRkJXVvlRHkpsKNQL<=0; 
			eKWoIeUrKiPbRIhuWEla<=0; 
			JRsyUSbxyBGBNdlJquOD<=0; 
			mobFFnIZQLEDGamGRCMQ<=0; 
			MIfRQTaujrTsVSIdukaO<=0; 
			qQxKziPkMaoHyxLiZQNv<=0; 
			SbGofGNBnFvEqTbzCMDT<=0; 
			eAyuUdQDmhsyVqUkrWtf<=0; 
			xcrfMbSpXdXRmlkuZRPx<=0; 
			BKSeIpcsVISDrrWyloru<=0; 
			cFxrUFXVhwbgFamPfIXu<=0; 
			EawSFufNSOZZHKtrbfDb<=0; 
			TtHHtKtzZHIcJuWziTSX<=0; 
			KAQFclKTjvNuQpWZONVn<=0; 
			zdDIxzPkCVYUHKycUMxS<=0; 
			yRWhBghWQtDlHOXzOKHV<=0; 
			xzEZrlRsvTQMlJcdcoBA<=0; 
			omKttYZtWwSNmJfXmNhw<=0; 
			TJsrTmKBrLuIryymjrla<=0; 
			UQIvtuLZLyNrLBcITiBh<=0; 
			dewJijMNQrULKORvfOPu<=0; 
			fFCHqQnaXGJtQcWhDHoo<=0; 
			lDVujeiDOsfmAcgTJEeH<=0; 
			tHYVLHNrDsWBBiksZJSh<=0; 
			YGcrryHhhucPWCRpoXpV<=0; 
			vhaFurczuHuVJndQizpm<=0; 
			bAUZnBUzAeFxTBCaAwBD<=0; 
			SJSSeEtWLefcHjjHknTt<=0; 
			RrXElmqzMleQDmHbRetu<=0; 
			RiwCfvabTaSgTyqQQkNP<=0; 
			ijLmWvKcGWYkfmVliDIH<=0; 
			JhZCVmRnYDVfDuTgaJBq<=0; 
			MmtedWLnvMwKkqgwBoYk<=0; 
			xNONPhZsuWCOqfHyKvVw<=0; 
			UYtsWPGzDLbsLPHFFzpM<=0; 
			HaIozTBrCuKZJRqUpAty<=0; 
			ihhBdoTzqImqsCjVxwKM<=0; 
			LPKCNZYNtyFJTUiKvFKI<=0; 
			VcDzTcOFndjUjhnRfxTN<=0; 
			ScSvdbbLcbwcpTKFudIt<=0; 
			ZFOGopcNcymIuYXsiiRw<=0; 
			zVAojGgdEwSIpPjTZZId<=0; 
			qwGWpRzKYsDLRvxcxAAH<=0; 
			WPkpODdzyINGGhuwZyoF<=0; 
			BaxiLnGgFxSKHVKkEWrL<=0; 
			cChsgcLGnvNEmegZREam<=0; 
			FRCWHcmIuMUUWgdYMzWu<=0; 
			QDYrIGBlnoXdNCUflHOP<=0; 
			zzYTnLgksIjwqZSweXMf<=0; 
			cWljGAlocPwsnrDyMjHO<=0; 
			JPYOnWGSGjFuHZfQBaEZ<=0; 
			VzfYJEwelHYPMpUSDmsC<=0; 
			XYQGKDohhXYVCeaCtmre<=0; 
			GbajCDnxXLGTStnsYsds<=0; 
			THlQvXwjkuLqdcMtPxBy<=0; 
			avkJIgYNFpvoyRkxaMTC<=0; 
			yhgnNUWIhVDlrtUDGEZn<=0; 
			lHvULbFfwhQgtqfjhwzH<=0; 
			TymwlUFeZUaLhFoWTZzU<=0; 
			obAWtmAwdFBYPXQlSuSy<=0; 
			VBJGcheVZYcxGpvcuBoi<=0; 
			NpcOSbiIpOcdgCjboENs<=0; 
			PiHYPPmDrZQNPnlqBFSt<=0; 
			rOXoAhCRFHntxISYSkye<=0; 
			IsXHeZVJKogNnFFfJwvx<=0; 
			BtfuDWbiQheMoNKySKtm<=0; 
			lsMUeaCgYLjCPUiUXaIc<=0; 
			kTdnGvNmLrhbepFdhZCh<=0; 
			vKbnovNlLRioZoJsQunL<=0; 
			nXBrtwwgIArkXUbHKAye<=0; 
			czvIYhYPaYPpRHUBJMFc<=0; 
			nsezjQWxmqwzmxCwosDv<=0; 
			ruIyZIesSthmxIaXEtrJ<=0; 
			cXQjLxPFTWRBhlJmdxUJ<=0; 
			GPoMmfciZsakCXuJMdbD<=0; 
			sZUCFycPxeatsZozmHJN<=0; 
			XbnmwpButuNSkogDlbQb<=0; 
			wdkDXnIkWnpQMmswGQeU<=0; 
			KpEHEcApUpQBvCLoAeYT<=0; 
			KsaghLmgaRvpRfCktbJZ<=0; 
			lZVGNfUlVmsuLbJxnQDA<=0; 
			rMBkqrLcKhflEMUYxGkE<=0; 
			wMlYFxkSbZTCTvhQOIei<=0; 
			WQGVbnQQZGQWVmpcxvbb<=0; 
			AzsKalhmBYUitbArLbcU<=0; 
			ekrMWzROxYoWtRpdbLZH<=0; 
			uLMmObkZiwzDlReqMwJN<=0; 
			eAEEsZkRTlfXOeEdICRO<=0; 
			DyXCiZssIzbywKGAbIwY<=0; 
			wBOVUPcFUWzhOUKDlJVa<=0; 
			BCsgCSHvysHWLteqbRMX<=0; 
			FrvVghZEElOfAJGPEURk<=0; 
			DHNpdfPdlvcIeMhPYCBD<=0; 
			ByKBiFClfZeeoBwNqVdH<=0; 
			muXlkjUrAqYazTUUGcVg<=0; 
			rZlIolWetZZffpSrlMAn<=0; 
			fCxfzzVrwjVhwiuAOpOD<=0; 
			VHDrEEGVFWccsKXzbEjD<=0; 
			pgbmZFwAnGMkExuHZexG<=0; 
			CYTIFZXRYHDOwAOpYhTY<=0; 
			hzujftnKaamrwjRBenpS<=0; 
			DwBiXGPwomcqrFUiwGKO<=0; 
			TxOTbaXnfvTWWAEMVKsT<=0; 
			VBPMSBgUzhZWqifRFXLt<=0; 
			fBEMznDkaUpJbucpUFUs<=0; 
			RXuUWWKfwotmzMaIdOHs<=0; 
			DScSrBltRCaJuMKRHxjp<=0; 
			yKhNJjIQvjuuxuKGtNvD<=0; 
			MBLbhXLxXGZHZERKIoYb<=0; 
			AiFthZhNPfZiXSnyPCOt<=0; 
			uDpYTElkHJsWMgegRIkv<=0; 
			LqJHECWMJlDdyFDTTZZH<=0; 
			ohfsyAOCKLVNdUfnlZGT<=0; 
			MOoDdDePAGBzQbLCZlwX<=0; 
			MHLazVdHgoSmGTltAxsJ<=0; 
			CYSqcBzpHDXSSATrgQjL<=0; 
			rPKZMoWgFDpDSJXXQmEU<=0; 
			hniufLGfdzmHbDIvsTIo<=0; 
			wTfPVycgpDcgGCOQhJjH<=0; 
			lcOMvsbHZmIJccXoDkqZ<=0; 
			UKirjTCurmcGUGGogrnh<=0; 
			KVLRCNcgwgdezgxdbtiz<=0; 
			ISUkQBFCDDhkmXDnEdVT<=0; 
			wLiUXxuAUdxCuAoAbUxH<=0; 
			vQNMUmgdbJJDFKzsjqLK<=0; 
			PPaVHoPQXNFqYDIgCroQ<=0; 
			fZmgOJpwMcdeRjEcecxZ<=0; 
			pXxRQDEgUJLwgwAsNvmV<=0; 
			JWyFVCrskBwarfgMzbIK<=0; 
			nLMIykvKsueQiebJRjaB<=0; 
			MwUAnLVNdEpwKFXarSrE<=0; 
			rwKFeNNlWzDutFvKudZd<=0; 
			YFTuhpacOohGrtlEUgyn<=0; 
			orsjfJIPQQvjIhvrnfZT<=0; 
			beooHOrejCcWcSXDuAMs<=0; 
			wLFqLqnhtGKyjhXVaXLu<=0; 
			VhlEwlgxfirfMpIAJZhE<=0; 
			ybSCwixJTEhXYyRpEeDj<=0; 
			PLAwknGzfcioZVaFOQCX<=0; 
			WdDdHRBJZdBPCxmYbWdk<=0; 
			BIxIzsQvWljjGYxMCQtS<=0; 
			TZYUrtPvAdyOAezlYVJO<=0; 
			qPqZhRZBobhmAXNGrsmh<=0; 
			BCGaGkllXBcyohBosHqS<=0; 
			pcgiabuotmBHXKOYDDAq<=0; 
			VidvAsXIfsppEpKtZeYc<=0; 
			lGfaCxQtDihDBzWEuyaH<=0; 
			ucwrtDfHQDZIjkmTmCvN<=0; 
			dayIzRpYaQRnEjXynbCm<=0; 
			vqgpItmCwuhiwKZyFXMt<=0; 
			FnVEwsGKlXZfUqxZGqHn<=0; 
			bitnzrgsExKEWSXnsRZq<=0; 
			eYsNwIgUOqnSppAZBKfW<=0; 
			FXTNpbkOJRifihZRkFUk<=0; 
			UCyPKegIVHgIqztViRHP<=0; 
			urwbynurHojveDuzQAqY<=0; 
			djsdiJHbeUEoOocTIVAL<=0; 
			juEeWiBDxjlSPOBoDWca<=0; 
			ZfhQiwfaJoKgwqVVBKhf<=0; 
			SNnVNrhdPUfxhixiespl<=0; 
			cHHoYqPSIzoxFEuXvNLY<=0; 
			hLpCUWbILJOjqbDhVEwn<=0; 
			itXQCyFacJzvPyzfGwVe<=0; 
			iujmIQQClXPYAKjueUBD<=0; 
			BjdcbpGuKPxnpZzFTfte<=0; 
			ZQFzyLJsVraTCGkqQcZA<=0; 
			fADZyEOwTyWvSQFgOnwG<=0; 
			xbhqvpXrDTlnyBNQeAlC<=0; 
			usigvHtlPqTHmByMEGLy<=0; 
			EqRnSoIxQaLPlCNmpBmq<=0; 
			VzsEzvUFwafgXDXiMnOI<=0; 
			qjQChEpAPSbKmoDGRppN<=0; 
			XBdmfGxuWrXGMBFOANKF<=0; 
			iHWmgCopJntOccGPObxn<=0; 
			eeoTbTyuwxPCsjuUGnLj<=0; 
			MkxrURKJtUzHVTfBwhoO<=0; 
			USFkaPtDBVOjbGpLXKUX<=0; 
			xcBSpPXNgyeMCKwBcsxX<=0; 
			APZhwjfiYOuKluWEaTIj<=0; 
			eiYeGwmYgODBCzcNuNtn<=0; 
			rmoQVcRSrSeskIibJzCc<=0; 
			AzSDmFqniQGEkrUvtcQd<=0; 
			BYQMYRDRDKXGHnLYQyKL<=0; 
			iYaojeeenaSObFkfIEyS<=0; 
			OvjWCALXGQonpSVNSUDx<=0; 
			QNSQONiKmlvpucXZsAKo<=0; 
			RKLbOFQSgMkwEdftvnBQ<=0; 
			hoPvrLDkwXFTkYESCUcp<=0; 
			hShwACbdYktXmGxyazAM<=0; 
			puehHutFkvCRvoGqbSYp<=0; 
			CSpvXCVkXjBnWvAFEiDG<=0; 
			GBnbMGmdJLNqPHpTRJqo<=0; 
			PQFlqUWXvhfFTKRniEDA<=0; 
			mNQfwTdWpUOnxIhbTYfU<=0; 
			ldQowZgtPeXlzjFcyWQl<=0; 
			HYWHYpKWyjTHzWIzGNeE<=0; 
			vsHmuANStIQsYgoNHsHw<=0; 
			tYWmIUymjXADFjUmKFpP<=0; 
			OQmggBTvOqhAXBiDJeaP<=0; 
			EFcUAERFHbivPwgHAMQa<=0; 
			jpbydIYGKyCwhjgemImi<=0; 
			OVYjPuZDVHOTTeuFPkrT<=0; 
			DqhwOfIUxBzsVSgEjWzC<=0; 
			plztNCDwyKBliboMvXKs<=0; 
			GojVETmCGfWcYwVYimBv<=0; 
			aogDiFiAXQqphSrsQbJV<=0; 
			rCOKgSoVLfXaUWFdsBnJ<=0; 
			ZuONZDcmHxALaUULMEAA<=0; 
			KIjEeYrBOSrzUMqGYBsV<=0; 
			ZBocacKljeyYorCiQgzQ<=0; 
			mqazMnBgYnlLqLRzaNYx<=0; 
			oyfKvpCwkpoCCxTglCJr<=0; 
			NGNEGckWnRLaqnjOKOmx<=0; 
			cVWqyzzrUUodYFbrorBz<=0; 
			RjwugczIYXEQzzmUrnYh<=0; 
			lEqWgKBWIbLvYwrXeDtN<=0; 
			DhnZhzYLzUMXzuxLMdpR<=0; 
			WwogGcAbNuwPRaXHfllR<=0; 
			fymbKnqnRYaHIRuPXxle<=0; 
			nJWkhXEkUmrasSyMThpL<=0; 
			qXNWBYTrrKKKGSroThrT<=0; 
			OWgmvdYcTEmvwkEuDkJS<=0; 
			urpaOisfjSiDXEZoTBsG<=0; 
			mveotDylkopgLZJFFBVl<=0; 
			CCXECvtOeIBEOFePtIRw<=0; 
			iYYwLjjGMjLikfxxrxIB<=0; 
			BJhcDugYXUoZuTXYBzJg<=0; 
			wpEZHrezpouBVvAiIOpn<=0; 
			omjfRcaEwaSdXWjgQYUv<=0; 
			aWXCrpICnOAsyXgkDTDT<=0; 
			HjXRkNnhDmrrYeoZLfga<=0; 
			zDWiKpAenkhcNZIBSNiT<=0; 
			UfyNbuBOwMXEdumKnlqN<=0; 
			LYSwVHbgNGVrAkuDLmxY<=0;
		end
		else if(gStNdqadtalDMswfRuqW==SHIFT_PASS_FIRST_HEADER)
		begin
			case(OhIQvlSNredlAvEzVwlD)                 
				1  :MNhKBwmQfBNRRoCGsGYL  <=MNhKBwmQfBNRRoCGsGYL  +CHmFHLXDhsSOMWPfgbXw;
				2  :CZUlnpSgUmTCmXxNawKq  <=CZUlnpSgUmTCmXxNawKq  +CHmFHLXDhsSOMWPfgbXw;
				3  :GCKDpTZdSkziHIHQTHTY  <=GCKDpTZdSkziHIHQTHTY  +CHmFHLXDhsSOMWPfgbXw;
				4  :TbggffYtMBhiLSACnOtm  <=TbggffYtMBhiLSACnOtm  +CHmFHLXDhsSOMWPfgbXw;
				5  :QMFreKPqLMtYHbzgqBQA  <=QMFreKPqLMtYHbzgqBQA  +CHmFHLXDhsSOMWPfgbXw;
				6  :NlcVQzrrHSpHBCrquBjt  <=NlcVQzrrHSpHBCrquBjt  +CHmFHLXDhsSOMWPfgbXw;
				7  :FSYqURbHbEaesQcTkdrx  <=FSYqURbHbEaesQcTkdrx  +CHmFHLXDhsSOMWPfgbXw;
				8  :qEtkygphCMCbDqrWtklY  <=qEtkygphCMCbDqrWtklY  +CHmFHLXDhsSOMWPfgbXw;
				9  :TLjaqwEsoHtrvWTBQRsK  <=TLjaqwEsoHtrvWTBQRsK  +CHmFHLXDhsSOMWPfgbXw;
				10 :cYsREsbuuQNtJwVuIQtc <=cYsREsbuuQNtJwVuIQtc +CHmFHLXDhsSOMWPfgbXw;
				11 :IADijSHmLDuBqTQJOxSa <=IADijSHmLDuBqTQJOxSa +CHmFHLXDhsSOMWPfgbXw;
				12 :BhAYLsocIYeStsZZVTUF <=BhAYLsocIYeStsZZVTUF +CHmFHLXDhsSOMWPfgbXw;
				13 :WQWSkTgEaMFMXPEsFHwg <=WQWSkTgEaMFMXPEsFHwg +CHmFHLXDhsSOMWPfgbXw;
				14 :WVikipTMfwFUtPMyACXK <=WVikipTMfwFUtPMyACXK +CHmFHLXDhsSOMWPfgbXw;
				15 :dXrKEPxqSBOppMxaytbW <=dXrKEPxqSBOppMxaytbW +CHmFHLXDhsSOMWPfgbXw;
				16 :NnjJwuwNoVWroSgcnSsE <=NnjJwuwNoVWroSgcnSsE +CHmFHLXDhsSOMWPfgbXw;
				17 :ASCWICejFoBbZHMJMVyD <=ASCWICejFoBbZHMJMVyD +CHmFHLXDhsSOMWPfgbXw;
				18 :twyoccXqjNTyiiCHZKgQ <=twyoccXqjNTyiiCHZKgQ +CHmFHLXDhsSOMWPfgbXw;
				19 :xvRCARkQSEXoZFEiGfjC <=xvRCARkQSEXoZFEiGfjC +CHmFHLXDhsSOMWPfgbXw;
				20 :JjLGddxBYbYmoYBVjdju <=JjLGddxBYbYmoYBVjdju +CHmFHLXDhsSOMWPfgbXw;
				21 :xyvvBnpUfpnejSAdOrIU <=xyvvBnpUfpnejSAdOrIU +CHmFHLXDhsSOMWPfgbXw;
				22 :LNWqJGCGvJkqDqnyFdST <=LNWqJGCGvJkqDqnyFdST +CHmFHLXDhsSOMWPfgbXw;
				23 :XXnujvRmwKtqZZbYXNom <=XXnujvRmwKtqZZbYXNom +CHmFHLXDhsSOMWPfgbXw;
				24 :rdgcYAhdMEGqsgkVVhHB <=rdgcYAhdMEGqsgkVVhHB +CHmFHLXDhsSOMWPfgbXw;
				25 :bcCzAdPYbGFOdbqFGtNY <=bcCzAdPYbGFOdbqFGtNY +CHmFHLXDhsSOMWPfgbXw;
				26 :MRTHuncHaQWNXrTdnjLu <=MRTHuncHaQWNXrTdnjLu +CHmFHLXDhsSOMWPfgbXw;
				27 :ZqxWPnvGQEisPGNSDkWt <=ZqxWPnvGQEisPGNSDkWt +CHmFHLXDhsSOMWPfgbXw;
				28 :jLboxjBIZGftrbnYaDHz <=jLboxjBIZGftrbnYaDHz +CHmFHLXDhsSOMWPfgbXw;
				29 :XPHrltKlkTYeddIYErlL <=XPHrltKlkTYeddIYErlL +CHmFHLXDhsSOMWPfgbXw;
				30 :DwnEuDbYEGceHCFfntWU <=DwnEuDbYEGceHCFfntWU +CHmFHLXDhsSOMWPfgbXw;
				31 :AhXRxsizDLdrPCSJbgvu <=AhXRxsizDLdrPCSJbgvu +CHmFHLXDhsSOMWPfgbXw;
				32 :dRLKJNMhCWjmYIXyBBMS <=dRLKJNMhCWjmYIXyBBMS +CHmFHLXDhsSOMWPfgbXw;
				33 :qKakmPsWXvxWDjopwmhd <=qKakmPsWXvxWDjopwmhd +CHmFHLXDhsSOMWPfgbXw;
				34 :OfKBQrlHgohHRFQMqPuX <=OfKBQrlHgohHRFQMqPuX +CHmFHLXDhsSOMWPfgbXw;
				35 :OMUVfbzXJtBmpgGUlWIN <=OMUVfbzXJtBmpgGUlWIN +CHmFHLXDhsSOMWPfgbXw;
				36 :pRjKNldSGgrOVpMtRdhl <=pRjKNldSGgrOVpMtRdhl +CHmFHLXDhsSOMWPfgbXw;
				37 :FzItXojZYuRrQPYroXqa <=FzItXojZYuRrQPYroXqa +CHmFHLXDhsSOMWPfgbXw;
				38 :tiASKMApdODRGubKCrIk <=tiASKMApdODRGubKCrIk +CHmFHLXDhsSOMWPfgbXw;
				39 :AofWIQWGCHGeAWxyBSnX <=AofWIQWGCHGeAWxyBSnX +CHmFHLXDhsSOMWPfgbXw;
				40 :BVZJHRZIRDJUNzlhOXNj <=BVZJHRZIRDJUNzlhOXNj +CHmFHLXDhsSOMWPfgbXw;
				41 :MJngMbRNrQAqZKOoJbfA <=MJngMbRNrQAqZKOoJbfA +CHmFHLXDhsSOMWPfgbXw;
				42 :LKEbaiUcnUkcdhTlxIWn <=LKEbaiUcnUkcdhTlxIWn +CHmFHLXDhsSOMWPfgbXw;
				43 :PIdKWDjIZqdVETXVKUyz <=PIdKWDjIZqdVETXVKUyz +CHmFHLXDhsSOMWPfgbXw;
				44 :TeweoifYlvYAXegPEOev <=TeweoifYlvYAXegPEOev +CHmFHLXDhsSOMWPfgbXw;
				45 :aHdPRBehEsBXhVSVEVGI <=aHdPRBehEsBXhVSVEVGI +CHmFHLXDhsSOMWPfgbXw;
				46 :EHDzFoGEUiKMcpmeZndO <=EHDzFoGEUiKMcpmeZndO +CHmFHLXDhsSOMWPfgbXw;
				47 :iGWdFxfLkcoPAfSnTRiW <=iGWdFxfLkcoPAfSnTRiW +CHmFHLXDhsSOMWPfgbXw;
				48 :OgwvxakMlGIDTjsTTTrF <=OgwvxakMlGIDTjsTTTrF +CHmFHLXDhsSOMWPfgbXw;
				49 :hweOwCSFFCFpnLABsNDz <=hweOwCSFFCFpnLABsNDz +CHmFHLXDhsSOMWPfgbXw;
				50 :kFILldZgHWqtwHcEyrEz <=kFILldZgHWqtwHcEyrEz +CHmFHLXDhsSOMWPfgbXw;
				51 :BHxWpRKaPloRmedcGnVS <=BHxWpRKaPloRmedcGnVS +CHmFHLXDhsSOMWPfgbXw;
				52 :jEDhTzjvJVSeQkYxJusx <=jEDhTzjvJVSeQkYxJusx +CHmFHLXDhsSOMWPfgbXw;
				53 :nVWwCingLJiAmNkXNBse <=nVWwCingLJiAmNkXNBse +CHmFHLXDhsSOMWPfgbXw;
				54 :hdQpCNCsCpWxWjyDHYIf <=hdQpCNCsCpWxWjyDHYIf +CHmFHLXDhsSOMWPfgbXw;
				55 :mYfjBwhqQaPjGDGuVzVT <=mYfjBwhqQaPjGDGuVzVT +CHmFHLXDhsSOMWPfgbXw;
				56 :sPdTjZhZROmcYPkfxnHK <=sPdTjZhZROmcYPkfxnHK +CHmFHLXDhsSOMWPfgbXw;
				57 :VOSkkJBkJQjLTSFCXXZG <=VOSkkJBkJQjLTSFCXXZG +CHmFHLXDhsSOMWPfgbXw;
				58 :wnDMhVWFcihAknOuJWgt <=wnDMhVWFcihAknOuJWgt +CHmFHLXDhsSOMWPfgbXw;
				59 :ZJYNMlOSJujZtBMVfIcG <=ZJYNMlOSJujZtBMVfIcG +CHmFHLXDhsSOMWPfgbXw;
				60 :cUQgUjrarAoCxWvadhrh <=cUQgUjrarAoCxWvadhrh +CHmFHLXDhsSOMWPfgbXw;
				61 :ayPBmMeTERtfSkylBBkl <=ayPBmMeTERtfSkylBBkl +CHmFHLXDhsSOMWPfgbXw;
				62 :zjiIArXGbkjgPxxXfPxg <=zjiIArXGbkjgPxxXfPxg +CHmFHLXDhsSOMWPfgbXw;
				63 :YERHnxdykgyyioNNZJSQ <=YERHnxdykgyyioNNZJSQ +CHmFHLXDhsSOMWPfgbXw;
				64 :rNuBwbgCniYGlSgOMCnE <=rNuBwbgCniYGlSgOMCnE +CHmFHLXDhsSOMWPfgbXw;
				65 :VjtVxkxLZrdVPkMsyEqe <=VjtVxkxLZrdVPkMsyEqe +CHmFHLXDhsSOMWPfgbXw;
				66 :fFwIafFNLTVTiIeJUZOi <=fFwIafFNLTVTiIeJUZOi +CHmFHLXDhsSOMWPfgbXw;
				67 :JofSpHHAILpRCvnGOmzf <=JofSpHHAILpRCvnGOmzf +CHmFHLXDhsSOMWPfgbXw;
				68 :OeYMhMfjeDdvkecHiLUT <=OeYMhMfjeDdvkecHiLUT +CHmFHLXDhsSOMWPfgbXw;
				69 :tVOTCptQSOpsjFBXiksw <=tVOTCptQSOpsjFBXiksw +CHmFHLXDhsSOMWPfgbXw;
				70 :AhXuWEaSPuUvIcwDuFWr <=AhXuWEaSPuUvIcwDuFWr +CHmFHLXDhsSOMWPfgbXw;
				71 :ekQuaIqPJyasZNSLaQOo <=ekQuaIqPJyasZNSLaQOo +CHmFHLXDhsSOMWPfgbXw;
				72 :osvtoSWcIuWcmvZruLsS <=osvtoSWcIuWcmvZruLsS +CHmFHLXDhsSOMWPfgbXw;
				73 :BzXYfwLRzqKLxtfxvmZC <=BzXYfwLRzqKLxtfxvmZC +CHmFHLXDhsSOMWPfgbXw;
				74 :tgVDzxwqtPquEcvdvFrC <=tgVDzxwqtPquEcvdvFrC +CHmFHLXDhsSOMWPfgbXw;
				75 :DzNsyDbNrzFrSyvQMHnd <=DzNsyDbNrzFrSyvQMHnd +CHmFHLXDhsSOMWPfgbXw;
				76 :iOnjZhBOoaDLaXXeVrwx <=iOnjZhBOoaDLaXXeVrwx +CHmFHLXDhsSOMWPfgbXw;
				77 :XwvNGtBVJXErWQRUuqBI <=XwvNGtBVJXErWQRUuqBI +CHmFHLXDhsSOMWPfgbXw;
				78 :JJgTPGsdUTcAdufkeJgK <=JJgTPGsdUTcAdufkeJgK +CHmFHLXDhsSOMWPfgbXw;
				79 :TfnRFMUqcGKfwYVkrOcp <=TfnRFMUqcGKfwYVkrOcp +CHmFHLXDhsSOMWPfgbXw;
				80 :kuHTqKTEGHJGjcgKEkCF <=kuHTqKTEGHJGjcgKEkCF +CHmFHLXDhsSOMWPfgbXw;
				81 :FfvTBiXNEwWARzrRMUYh <=FfvTBiXNEwWARzrRMUYh +CHmFHLXDhsSOMWPfgbXw;
				82 :VMfdRrsDolDymeMDbscN <=VMfdRrsDolDymeMDbscN +CHmFHLXDhsSOMWPfgbXw;
				83 :iPuXoTiWLBGZVYAHGaYO <=iPuXoTiWLBGZVYAHGaYO +CHmFHLXDhsSOMWPfgbXw;
				84 :BaxkmTikPlEanrOALJQn <=BaxkmTikPlEanrOALJQn +CHmFHLXDhsSOMWPfgbXw;
				85 :TGPYgdsEOqsHqlpqyhVp <=TGPYgdsEOqsHqlpqyhVp +CHmFHLXDhsSOMWPfgbXw;
				86 :VZaWDekOPjcbcuLkmTCK <=VZaWDekOPjcbcuLkmTCK +CHmFHLXDhsSOMWPfgbXw;
				87 :ceSSpUnFGIqusvzAQYyv <=ceSSpUnFGIqusvzAQYyv +CHmFHLXDhsSOMWPfgbXw;
				88 :KkgZHqKRoBphLNurbXZv <=KkgZHqKRoBphLNurbXZv +CHmFHLXDhsSOMWPfgbXw;
				89 :BVfKHJmimWhfvhFZYdJC <=BVfKHJmimWhfvhFZYdJC +CHmFHLXDhsSOMWPfgbXw;
				90 :XWIoNGOmiUqZuWDNerJA <=XWIoNGOmiUqZuWDNerJA +CHmFHLXDhsSOMWPfgbXw;
				91 :ymZNoaOSvkuMNFrKCZJc <=ymZNoaOSvkuMNFrKCZJc +CHmFHLXDhsSOMWPfgbXw;
				92 :JtPboWbpZfxqTBEEDYyf <=JtPboWbpZfxqTBEEDYyf +CHmFHLXDhsSOMWPfgbXw;
				93 :NIzOkTmOrsmtdJpYgwkn <=NIzOkTmOrsmtdJpYgwkn +CHmFHLXDhsSOMWPfgbXw;
				94 :HPBVjcjYzqThfAZsuBko <=HPBVjcjYzqThfAZsuBko +CHmFHLXDhsSOMWPfgbXw;
				95 :RtOUSNvLjifycdHERnsH <=RtOUSNvLjifycdHERnsH +CHmFHLXDhsSOMWPfgbXw;
				96 :RHqjRVMUmlsTYhhiTxqt <=RHqjRVMUmlsTYhhiTxqt +CHmFHLXDhsSOMWPfgbXw;
				97 :irQWRPjnSymTgyEWfOeV <=irQWRPjnSymTgyEWfOeV +CHmFHLXDhsSOMWPfgbXw;
				98 :gHMMxJFDpgQtSoSKsfzc <=gHMMxJFDpgQtSoSKsfzc +CHmFHLXDhsSOMWPfgbXw;
				99 :XrXzzUeQwqtdbHighLXh <=XrXzzUeQwqtdbHighLXh +CHmFHLXDhsSOMWPfgbXw;
				100:VXesUOJyNaYiksaASUmr<=VXesUOJyNaYiksaASUmr+CHmFHLXDhsSOMWPfgbXw; 
				101:MjDYzSbWZYtgtBPeFxFX<=MjDYzSbWZYtgtBPeFxFX+CHmFHLXDhsSOMWPfgbXw; 
				102:QocIghyhzPXBoGjaFxEW<=QocIghyhzPXBoGjaFxEW+CHmFHLXDhsSOMWPfgbXw; 
				103:aNNRDAQndlQbuwTNoeBC<=aNNRDAQndlQbuwTNoeBC+CHmFHLXDhsSOMWPfgbXw; 
				104:ganwYnOuHsVFGlnGQGGf<=ganwYnOuHsVFGlnGQGGf+CHmFHLXDhsSOMWPfgbXw; 
				105:TmUIbPULspEIyexiGCHU<=TmUIbPULspEIyexiGCHU+CHmFHLXDhsSOMWPfgbXw; 
				106:GrWFHsoruHLBTofZiNlc<=GrWFHsoruHLBTofZiNlc+CHmFHLXDhsSOMWPfgbXw; 
				107:HemnvXRItkGWOQQBARSS<=HemnvXRItkGWOQQBARSS+CHmFHLXDhsSOMWPfgbXw; 
				108:crDvxwhExTyEkehZAJBR<=crDvxwhExTyEkehZAJBR+CHmFHLXDhsSOMWPfgbXw; 
				109:vqFRiEdZYIvaYIjwIZPo<=vqFRiEdZYIvaYIjwIZPo+CHmFHLXDhsSOMWPfgbXw; 
				110:RiyBtzLqNImqdjYXxYLF<=RiyBtzLqNImqdjYXxYLF+CHmFHLXDhsSOMWPfgbXw; 
				111:QAZelRxmduKrKymXyprg<=QAZelRxmduKrKymXyprg+CHmFHLXDhsSOMWPfgbXw; 
				112:IixlIEeyecDFQCcIcXFK<=IixlIEeyecDFQCcIcXFK+CHmFHLXDhsSOMWPfgbXw; 
				113:CahtEzYLkeeOsdRKBvoI<=CahtEzYLkeeOsdRKBvoI+CHmFHLXDhsSOMWPfgbXw; 
				114:hXvwCaJPKLmTlGnIqShO<=hXvwCaJPKLmTlGnIqShO+CHmFHLXDhsSOMWPfgbXw; 
				115:ZapMeflJnJGQFrDdnzZx<=ZapMeflJnJGQFrDdnzZx+CHmFHLXDhsSOMWPfgbXw; 
				116:tEZVPsZbWePhmBDkYbkW<=tEZVPsZbWePhmBDkYbkW+CHmFHLXDhsSOMWPfgbXw; 
				117:VKIhSekuVtyFcvuoBpZH<=VKIhSekuVtyFcvuoBpZH+CHmFHLXDhsSOMWPfgbXw; 
				118:HHissIgZPvjjCfGzZWgP<=HHissIgZPvjjCfGzZWgP+CHmFHLXDhsSOMWPfgbXw; 
				119:ZthEdVQnyODdQJpzqpDX<=ZthEdVQnyODdQJpzqpDX+CHmFHLXDhsSOMWPfgbXw; 
				120:ZvVAYFyMKYuJjjuLlssM<=ZvVAYFyMKYuJjjuLlssM+CHmFHLXDhsSOMWPfgbXw; 
				121:BDVfxjBZqdgfpcXaqSxS<=BDVfxjBZqdgfpcXaqSxS+CHmFHLXDhsSOMWPfgbXw; 
				122:SYPrSAmIZhepjzRpfAbW<=SYPrSAmIZhepjzRpfAbW+CHmFHLXDhsSOMWPfgbXw; 
				123:bheecNbLIfuKFYksBrvM<=bheecNbLIfuKFYksBrvM+CHmFHLXDhsSOMWPfgbXw; 
				124:LoFfmBmHEBmQlYvRihJx<=LoFfmBmHEBmQlYvRihJx+CHmFHLXDhsSOMWPfgbXw; 
				125:RAqkMVQdcCkZqHQrYhTY<=RAqkMVQdcCkZqHQrYhTY+CHmFHLXDhsSOMWPfgbXw; 
				126:JwazcQrhGdLokRSxMIPy<=JwazcQrhGdLokRSxMIPy+CHmFHLXDhsSOMWPfgbXw; 
				127:NHwKTvStgXGxecepjZCb<=NHwKTvStgXGxecepjZCb+CHmFHLXDhsSOMWPfgbXw; 
				128:iFhOAEkrfnWgTHHMCrAr<=iFhOAEkrfnWgTHHMCrAr+CHmFHLXDhsSOMWPfgbXw; 
				129:KoZvZIhKhWDYlgwhYWfH<=KoZvZIhKhWDYlgwhYWfH+CHmFHLXDhsSOMWPfgbXw; 
				130:xqkVQlUmzixmBBOWsogM<=xqkVQlUmzixmBBOWsogM+CHmFHLXDhsSOMWPfgbXw; 
				131:mZcXpTwcGpwcsXaAXzJZ<=mZcXpTwcGpwcsXaAXzJZ+CHmFHLXDhsSOMWPfgbXw; 
				132:tBkJHywSnDHjCloeCKQN<=tBkJHywSnDHjCloeCKQN+CHmFHLXDhsSOMWPfgbXw; 
				133:rtIOwgMybhKPbMtTkPHH<=rtIOwgMybhKPbMtTkPHH+CHmFHLXDhsSOMWPfgbXw; 
				134:ULvOWCBpLiqodnUiPZne<=ULvOWCBpLiqodnUiPZne+CHmFHLXDhsSOMWPfgbXw; 
				135:UeCtXzcgpZHmscgLWNgU<=UeCtXzcgpZHmscgLWNgU+CHmFHLXDhsSOMWPfgbXw; 
				136:NchYslfTwDoJDaIhKQld<=NchYslfTwDoJDaIhKQld+CHmFHLXDhsSOMWPfgbXw; 
				137:vdLrgmXBDTPmGWwCZgJK<=vdLrgmXBDTPmGWwCZgJK+CHmFHLXDhsSOMWPfgbXw; 
				138:fypmfZbmWDbDCXEismjU<=fypmfZbmWDbDCXEismjU+CHmFHLXDhsSOMWPfgbXw; 
				139:FEgAuSjALENQXZOiGFUZ<=FEgAuSjALENQXZOiGFUZ+CHmFHLXDhsSOMWPfgbXw; 
				140:hUaTrhFAshrngFoHaXaJ<=hUaTrhFAshrngFoHaXaJ+CHmFHLXDhsSOMWPfgbXw; 
				141:avmhenqBbGIfSBAIabaF<=avmhenqBbGIfSBAIabaF+CHmFHLXDhsSOMWPfgbXw; 
				142:IlmCWYrxdJVqIQywKmAF<=IlmCWYrxdJVqIQywKmAF+CHmFHLXDhsSOMWPfgbXw; 
				143:GXKZdRvGRyUFWKyHVAFD<=GXKZdRvGRyUFWKyHVAFD+CHmFHLXDhsSOMWPfgbXw; 
				144:PExEfPxznaZHuROUSmfc<=PExEfPxznaZHuROUSmfc+CHmFHLXDhsSOMWPfgbXw; 
				145:DoWtmJCIdGMmwEInsyhi<=DoWtmJCIdGMmwEInsyhi+CHmFHLXDhsSOMWPfgbXw; 
				146:AtkWXjDVDEZLaumbWZzI<=AtkWXjDVDEZLaumbWZzI+CHmFHLXDhsSOMWPfgbXw; 
				147:HvOvrGAvaPTzYsRxiQFa<=HvOvrGAvaPTzYsRxiQFa+CHmFHLXDhsSOMWPfgbXw; 
				148:rwPuhbqaLGfEsTZJaDhF<=rwPuhbqaLGfEsTZJaDhF+CHmFHLXDhsSOMWPfgbXw; 
				149:YphfuswJNWiAbvgWEfjm<=YphfuswJNWiAbvgWEfjm+CHmFHLXDhsSOMWPfgbXw; 
				150:YhTJCIYfjiXccwQDAncB<=YhTJCIYfjiXccwQDAncB+CHmFHLXDhsSOMWPfgbXw; 
				151:KaDxyGuuayhqIxIwbGQG<=KaDxyGuuayhqIxIwbGQG+CHmFHLXDhsSOMWPfgbXw; 
				152:SCcERabQMmiRZhSuKFqS<=SCcERabQMmiRZhSuKFqS+CHmFHLXDhsSOMWPfgbXw; 
				153:ASVDnraQDtLQhInOEyVK<=ASVDnraQDtLQhInOEyVK+CHmFHLXDhsSOMWPfgbXw; 
				154:RzDedJWchbeEickgtFOM<=RzDedJWchbeEickgtFOM+CHmFHLXDhsSOMWPfgbXw; 
				155:qBWQIFhDbnPbANWZJPUR<=qBWQIFhDbnPbANWZJPUR+CHmFHLXDhsSOMWPfgbXw; 
				156:ONSywhEkLUpjhsBVzOEr<=ONSywhEkLUpjhsBVzOEr+CHmFHLXDhsSOMWPfgbXw; 
				157:SiWXyZwStCTfnlFxLPQx<=SiWXyZwStCTfnlFxLPQx+CHmFHLXDhsSOMWPfgbXw; 
				158:ljlzMOdncFtIKCHtOsVQ<=ljlzMOdncFtIKCHtOsVQ+CHmFHLXDhsSOMWPfgbXw; 
				159:sBtkXBZAHFHDVqMZHZdd<=sBtkXBZAHFHDVqMZHZdd+CHmFHLXDhsSOMWPfgbXw; 
				160:ZNywgghYzvszBznGurzE<=ZNywgghYzvszBznGurzE+CHmFHLXDhsSOMWPfgbXw; 
				161:giByCXZhzRJrKpUfJiYx<=giByCXZhzRJrKpUfJiYx+CHmFHLXDhsSOMWPfgbXw; 
				162:NOzoIRcSVgyFREyzzHqs<=NOzoIRcSVgyFREyzzHqs+CHmFHLXDhsSOMWPfgbXw; 
				163:hvcttLppSPcVixtVRHqN<=hvcttLppSPcVixtVRHqN+CHmFHLXDhsSOMWPfgbXw; 
				164:NXURaWZymtMESRzASoml<=NXURaWZymtMESRzASoml+CHmFHLXDhsSOMWPfgbXw; 
				165:OGJwXjhBDuVzMrVxGthI<=OGJwXjhBDuVzMrVxGthI+CHmFHLXDhsSOMWPfgbXw; 
				166:tDHSWWPwhDHPIdkjEtEW<=tDHSWWPwhDHPIdkjEtEW+CHmFHLXDhsSOMWPfgbXw; 
				167:spPgPLHCbVgdzOmJFakw<=spPgPLHCbVgdzOmJFakw+CHmFHLXDhsSOMWPfgbXw; 
				168:NCLfdSDEGhGvIWQaIuMS<=NCLfdSDEGhGvIWQaIuMS+CHmFHLXDhsSOMWPfgbXw; 
				169:NfdfbTCtNjYFDeLLecMe<=NfdfbTCtNjYFDeLLecMe+CHmFHLXDhsSOMWPfgbXw; 
				170:xIHGyzqgFJSHmjAJEkTk<=xIHGyzqgFJSHmjAJEkTk+CHmFHLXDhsSOMWPfgbXw; 
				171:ffdnbvLvbNGfaiXRKcYD<=ffdnbvLvbNGfaiXRKcYD+CHmFHLXDhsSOMWPfgbXw; 
				172:dDkKlvBKHVNSwGZicnzg<=dDkKlvBKHVNSwGZicnzg+CHmFHLXDhsSOMWPfgbXw; 
				173:sTYRbAXFBXVNlExKcFRO<=sTYRbAXFBXVNlExKcFRO+CHmFHLXDhsSOMWPfgbXw; 
				174:QYcegkQFzbKFzvlPxGeR<=QYcegkQFzbKFzvlPxGeR+CHmFHLXDhsSOMWPfgbXw; 
				175:WCbGOTtDaZUdMPlupDBN<=WCbGOTtDaZUdMPlupDBN+CHmFHLXDhsSOMWPfgbXw; 
				176:kNoeoxFOMGDTBbVzHlLM<=kNoeoxFOMGDTBbVzHlLM+CHmFHLXDhsSOMWPfgbXw; 
				177:pcsafTpJQiyaKivHSiiO<=pcsafTpJQiyaKivHSiiO+CHmFHLXDhsSOMWPfgbXw; 
				178:HhgKJaIdyWwhlApPzTKC<=HhgKJaIdyWwhlApPzTKC+CHmFHLXDhsSOMWPfgbXw; 
				179:LgxgHDHmFYbeGgXVWgvC<=LgxgHDHmFYbeGgXVWgvC+CHmFHLXDhsSOMWPfgbXw; 
				180:cKBOWdNoOXhznBHdAwlu<=cKBOWdNoOXhznBHdAwlu+CHmFHLXDhsSOMWPfgbXw; 
				181:KASZraJCWhbAUtfwnLfk<=KASZraJCWhbAUtfwnLfk+CHmFHLXDhsSOMWPfgbXw; 
				182:AGPbOkqoDAYNiAUBxYWb<=AGPbOkqoDAYNiAUBxYWb+CHmFHLXDhsSOMWPfgbXw; 
				183:QePGiiHhRVKoAUkzEcSD<=QePGiiHhRVKoAUkzEcSD+CHmFHLXDhsSOMWPfgbXw; 
				184:ULkqQHcjawmJPPtzcPCS<=ULkqQHcjawmJPPtzcPCS+CHmFHLXDhsSOMWPfgbXw; 
				185:gVMkJmsMEYFtEfiuwaKj<=gVMkJmsMEYFtEfiuwaKj+CHmFHLXDhsSOMWPfgbXw; 
				186:yHFGaozymIVZZMqtzLDd<=yHFGaozymIVZZMqtzLDd+CHmFHLXDhsSOMWPfgbXw; 
				187:XyhfMHNDiNoQgejMGALx<=XyhfMHNDiNoQgejMGALx+CHmFHLXDhsSOMWPfgbXw; 
				188:zWhpxSLccsmBmQBUhbQT<=zWhpxSLccsmBmQBUhbQT+CHmFHLXDhsSOMWPfgbXw; 
				189:xKWgakKpWyTQyBrwYCIS<=xKWgakKpWyTQyBrwYCIS+CHmFHLXDhsSOMWPfgbXw; 
				190:UkOdSdYxtcxumOakhLgx<=UkOdSdYxtcxumOakhLgx+CHmFHLXDhsSOMWPfgbXw; 
				191:nhnBLnxptnOVgbmRStCU<=nhnBLnxptnOVgbmRStCU+CHmFHLXDhsSOMWPfgbXw; 
				192:UmXpnIjWZNlfEPEYcDTn<=UmXpnIjWZNlfEPEYcDTn+CHmFHLXDhsSOMWPfgbXw; 
				193:deblhPqNAplcidEXSGqw<=deblhPqNAplcidEXSGqw+CHmFHLXDhsSOMWPfgbXw; 
				194:GgkZJHLDkhyFsCCzuqLa<=GgkZJHLDkhyFsCCzuqLa+CHmFHLXDhsSOMWPfgbXw; 
				195:pKDUrDrLLWTOdoUxvsyF<=pKDUrDrLLWTOdoUxvsyF+CHmFHLXDhsSOMWPfgbXw; 
				196:JrQYFpYwpBTANpnTvLiU<=JrQYFpYwpBTANpnTvLiU+CHmFHLXDhsSOMWPfgbXw; 
				197:KencLjTnnSFqjwbVxqJg<=KencLjTnnSFqjwbVxqJg+CHmFHLXDhsSOMWPfgbXw; 
				198:TXuaPuUIuhCkLiMhEKiF<=TXuaPuUIuhCkLiMhEKiF+CHmFHLXDhsSOMWPfgbXw; 
				199:aAhmLslHTfVKwKSRWVtp<=aAhmLslHTfVKwKSRWVtp+CHmFHLXDhsSOMWPfgbXw; 
				200:NJEYMnPHSmEVDftsqzQE<=NJEYMnPHSmEVDftsqzQE+CHmFHLXDhsSOMWPfgbXw; 
				201:ByBgtRovBsKUVHUQEzwk<=ByBgtRovBsKUVHUQEzwk+CHmFHLXDhsSOMWPfgbXw; 
				202:pcCSuYOgcgRTEfyKANVf<=pcCSuYOgcgRTEfyKANVf+CHmFHLXDhsSOMWPfgbXw; 
				203:OOJGXLeAUSSWDwWKvqMN<=OOJGXLeAUSSWDwWKvqMN+CHmFHLXDhsSOMWPfgbXw; 
				204:xzObOtBnVrtyMpWImLGp<=xzObOtBnVrtyMpWImLGp+CHmFHLXDhsSOMWPfgbXw; 
				205:fPvbFzCudNRdKXFIwPTW<=fPvbFzCudNRdKXFIwPTW+CHmFHLXDhsSOMWPfgbXw; 
				206:UCBlEpPTGRkqheRhrmew<=UCBlEpPTGRkqheRhrmew+CHmFHLXDhsSOMWPfgbXw; 
				207:rxGiYeZlkdsRNUfrmDKO<=rxGiYeZlkdsRNUfrmDKO+CHmFHLXDhsSOMWPfgbXw; 
				208:BRDRPJjxjaVvUmeEcabW<=BRDRPJjxjaVvUmeEcabW+CHmFHLXDhsSOMWPfgbXw; 
				209:twevQhSVcRXlOWMZGHZH<=twevQhSVcRXlOWMZGHZH+CHmFHLXDhsSOMWPfgbXw; 
				210:hsPTsFDtcTjmyeddHGwC<=hsPTsFDtcTjmyeddHGwC+CHmFHLXDhsSOMWPfgbXw; 
				211:SnXYHdlnJsKNjOCDlAdk<=SnXYHdlnJsKNjOCDlAdk+CHmFHLXDhsSOMWPfgbXw; 
				212:fzPjNCWXNlBXDEixcMfx<=fzPjNCWXNlBXDEixcMfx+CHmFHLXDhsSOMWPfgbXw; 
				213:MzxTqhCibhKKovZUinvJ<=MzxTqhCibhKKovZUinvJ+CHmFHLXDhsSOMWPfgbXw; 
				214:UjBCIuRFDGUvCwBBwjtv<=UjBCIuRFDGUvCwBBwjtv+CHmFHLXDhsSOMWPfgbXw; 
				215:WLvkMHkFFjSeXeCMFLqU<=WLvkMHkFFjSeXeCMFLqU+CHmFHLXDhsSOMWPfgbXw; 
				216:OdXRCGgZgKmtknFfVeGS<=OdXRCGgZgKmtknFfVeGS+CHmFHLXDhsSOMWPfgbXw; 
				217:YTagschVaYsVmCoZyGxw<=YTagschVaYsVmCoZyGxw+CHmFHLXDhsSOMWPfgbXw; 
				218:uBDeqwBeWjkFnJPifZac<=uBDeqwBeWjkFnJPifZac+CHmFHLXDhsSOMWPfgbXw; 
				219:ChqdVbAPIMvlcdCLZFDM<=ChqdVbAPIMvlcdCLZFDM+CHmFHLXDhsSOMWPfgbXw; 
				220:xVhIWQmsjbKYhycXOZZj<=xVhIWQmsjbKYhycXOZZj+CHmFHLXDhsSOMWPfgbXw; 
				221:moXSbLoysxSoGKFutzbo<=moXSbLoysxSoGKFutzbo+CHmFHLXDhsSOMWPfgbXw; 
				222:pFrrbOJSlADGwICgxTdA<=pFrrbOJSlADGwICgxTdA+CHmFHLXDhsSOMWPfgbXw; 
				223:eFKOOLSSWbJGsojVvoDI<=eFKOOLSSWbJGsojVvoDI+CHmFHLXDhsSOMWPfgbXw; 
				224:CjkyDsWsnyjeHKnTfjoz<=CjkyDsWsnyjeHKnTfjoz+CHmFHLXDhsSOMWPfgbXw; 
				225:ikgPtqNHSxOonFiPgvOK<=ikgPtqNHSxOonFiPgvOK+CHmFHLXDhsSOMWPfgbXw; 
				226:JzYgxPBzYqfsNCHdKwWT<=JzYgxPBzYqfsNCHdKwWT+CHmFHLXDhsSOMWPfgbXw; 
				227:rYlFPAhuURCPKCloqLOG<=rYlFPAhuURCPKCloqLOG+CHmFHLXDhsSOMWPfgbXw; 
				228:PQEjeJZSeiJdTNkqSiiS<=PQEjeJZSeiJdTNkqSiiS+CHmFHLXDhsSOMWPfgbXw; 
				229:MSaMrnCOKHvvWjrvrLVh<=MSaMrnCOKHvvWjrvrLVh+CHmFHLXDhsSOMWPfgbXw; 
				230:bZovfeygdcHHRKfkxfHl<=bZovfeygdcHHRKfkxfHl+CHmFHLXDhsSOMWPfgbXw; 
				231:ATkQsyvByLEkPXEmCGoF<=ATkQsyvByLEkPXEmCGoF+CHmFHLXDhsSOMWPfgbXw; 
				232:uBtJXFukNYPqTHWppmdv<=uBtJXFukNYPqTHWppmdv+CHmFHLXDhsSOMWPfgbXw; 
				233:soNzOmONAzHkpLFWdCtg<=soNzOmONAzHkpLFWdCtg+CHmFHLXDhsSOMWPfgbXw; 
				234:lLJeyDbtTaFvkSfqLcWK<=lLJeyDbtTaFvkSfqLcWK+CHmFHLXDhsSOMWPfgbXw; 
				235:lMFLPXTVXadwnVsRrAPI<=lMFLPXTVXadwnVsRrAPI+CHmFHLXDhsSOMWPfgbXw; 
				236:WPsXEglrQBPoHLKokyap<=WPsXEglrQBPoHLKokyap+CHmFHLXDhsSOMWPfgbXw; 
				237:RqjRxpMaojbkWLGINNMj<=RqjRxpMaojbkWLGINNMj+CHmFHLXDhsSOMWPfgbXw; 
				238:CcpgUvVvfmeEoXXGYlgz<=CcpgUvVvfmeEoXXGYlgz+CHmFHLXDhsSOMWPfgbXw; 
				239:yNeJpDTKbQScFfOFsIMP<=yNeJpDTKbQScFfOFsIMP+CHmFHLXDhsSOMWPfgbXw; 
				240:uVWYpFOIjqHtdFWqJLJL<=uVWYpFOIjqHtdFWqJLJL+CHmFHLXDhsSOMWPfgbXw; 
				241:vCLJZIRyvOOZpamupbmS<=vCLJZIRyvOOZpamupbmS+CHmFHLXDhsSOMWPfgbXw; 
				242:JiRCGeWXVDSjvohYatoO<=JiRCGeWXVDSjvohYatoO+CHmFHLXDhsSOMWPfgbXw; 
				243:JXVeYnVHSdAGpxmDHgjf<=JXVeYnVHSdAGpxmDHgjf+CHmFHLXDhsSOMWPfgbXw; 
				244:iXlLoGyimBUgUkjZoGvT<=iXlLoGyimBUgUkjZoGvT+CHmFHLXDhsSOMWPfgbXw; 
				245:JrBVZVJGLbQlQIuxVRMO<=JrBVZVJGLbQlQIuxVRMO+CHmFHLXDhsSOMWPfgbXw; 
				246:MZLrRshlRErhPsqJeccP<=MZLrRshlRErhPsqJeccP+CHmFHLXDhsSOMWPfgbXw; 
				247:KddqRkJXVvlRHkpsKNQL<=KddqRkJXVvlRHkpsKNQL+CHmFHLXDhsSOMWPfgbXw; 
				248:eKWoIeUrKiPbRIhuWEla<=eKWoIeUrKiPbRIhuWEla+CHmFHLXDhsSOMWPfgbXw; 
				249:JRsyUSbxyBGBNdlJquOD<=JRsyUSbxyBGBNdlJquOD+CHmFHLXDhsSOMWPfgbXw; 
				250:mobFFnIZQLEDGamGRCMQ<=mobFFnIZQLEDGamGRCMQ+CHmFHLXDhsSOMWPfgbXw; 
				251:MIfRQTaujrTsVSIdukaO<=MIfRQTaujrTsVSIdukaO+CHmFHLXDhsSOMWPfgbXw; 
				252:qQxKziPkMaoHyxLiZQNv<=qQxKziPkMaoHyxLiZQNv+CHmFHLXDhsSOMWPfgbXw; 
				253:SbGofGNBnFvEqTbzCMDT<=SbGofGNBnFvEqTbzCMDT+CHmFHLXDhsSOMWPfgbXw; 
				254:eAyuUdQDmhsyVqUkrWtf<=eAyuUdQDmhsyVqUkrWtf+CHmFHLXDhsSOMWPfgbXw; 
				255:xcrfMbSpXdXRmlkuZRPx<=xcrfMbSpXdXRmlkuZRPx+CHmFHLXDhsSOMWPfgbXw; 
				256:BKSeIpcsVISDrrWyloru<=BKSeIpcsVISDrrWyloru+CHmFHLXDhsSOMWPfgbXw; 
				257:cFxrUFXVhwbgFamPfIXu<=cFxrUFXVhwbgFamPfIXu+CHmFHLXDhsSOMWPfgbXw; 
				258:EawSFufNSOZZHKtrbfDb<=EawSFufNSOZZHKtrbfDb+CHmFHLXDhsSOMWPfgbXw; 
				259:TtHHtKtzZHIcJuWziTSX<=TtHHtKtzZHIcJuWziTSX+CHmFHLXDhsSOMWPfgbXw; 
				260:KAQFclKTjvNuQpWZONVn<=KAQFclKTjvNuQpWZONVn+CHmFHLXDhsSOMWPfgbXw; 
				261:zdDIxzPkCVYUHKycUMxS<=zdDIxzPkCVYUHKycUMxS+CHmFHLXDhsSOMWPfgbXw; 
				262:yRWhBghWQtDlHOXzOKHV<=yRWhBghWQtDlHOXzOKHV+CHmFHLXDhsSOMWPfgbXw; 
				263:xzEZrlRsvTQMlJcdcoBA<=xzEZrlRsvTQMlJcdcoBA+CHmFHLXDhsSOMWPfgbXw; 
				264:omKttYZtWwSNmJfXmNhw<=omKttYZtWwSNmJfXmNhw+CHmFHLXDhsSOMWPfgbXw; 
				265:TJsrTmKBrLuIryymjrla<=TJsrTmKBrLuIryymjrla+CHmFHLXDhsSOMWPfgbXw; 
				266:UQIvtuLZLyNrLBcITiBh<=UQIvtuLZLyNrLBcITiBh+CHmFHLXDhsSOMWPfgbXw; 
				267:dewJijMNQrULKORvfOPu<=dewJijMNQrULKORvfOPu+CHmFHLXDhsSOMWPfgbXw; 
				268:fFCHqQnaXGJtQcWhDHoo<=fFCHqQnaXGJtQcWhDHoo+CHmFHLXDhsSOMWPfgbXw; 
				269:lDVujeiDOsfmAcgTJEeH<=lDVujeiDOsfmAcgTJEeH+CHmFHLXDhsSOMWPfgbXw; 
				270:tHYVLHNrDsWBBiksZJSh<=tHYVLHNrDsWBBiksZJSh+CHmFHLXDhsSOMWPfgbXw; 
				271:YGcrryHhhucPWCRpoXpV<=YGcrryHhhucPWCRpoXpV+CHmFHLXDhsSOMWPfgbXw; 
				272:vhaFurczuHuVJndQizpm<=vhaFurczuHuVJndQizpm+CHmFHLXDhsSOMWPfgbXw; 
				273:bAUZnBUzAeFxTBCaAwBD<=bAUZnBUzAeFxTBCaAwBD+CHmFHLXDhsSOMWPfgbXw; 
				274:SJSSeEtWLefcHjjHknTt<=SJSSeEtWLefcHjjHknTt+CHmFHLXDhsSOMWPfgbXw; 
				275:RrXElmqzMleQDmHbRetu<=RrXElmqzMleQDmHbRetu+CHmFHLXDhsSOMWPfgbXw; 
				276:RiwCfvabTaSgTyqQQkNP<=RiwCfvabTaSgTyqQQkNP+CHmFHLXDhsSOMWPfgbXw; 
				277:ijLmWvKcGWYkfmVliDIH<=ijLmWvKcGWYkfmVliDIH+CHmFHLXDhsSOMWPfgbXw; 
				278:JhZCVmRnYDVfDuTgaJBq<=JhZCVmRnYDVfDuTgaJBq+CHmFHLXDhsSOMWPfgbXw; 
				279:MmtedWLnvMwKkqgwBoYk<=MmtedWLnvMwKkqgwBoYk+CHmFHLXDhsSOMWPfgbXw; 
				280:xNONPhZsuWCOqfHyKvVw<=xNONPhZsuWCOqfHyKvVw+CHmFHLXDhsSOMWPfgbXw; 
				281:UYtsWPGzDLbsLPHFFzpM<=UYtsWPGzDLbsLPHFFzpM+CHmFHLXDhsSOMWPfgbXw; 
				282:HaIozTBrCuKZJRqUpAty<=HaIozTBrCuKZJRqUpAty+CHmFHLXDhsSOMWPfgbXw; 
				283:ihhBdoTzqImqsCjVxwKM<=ihhBdoTzqImqsCjVxwKM+CHmFHLXDhsSOMWPfgbXw; 
				284:LPKCNZYNtyFJTUiKvFKI<=LPKCNZYNtyFJTUiKvFKI+CHmFHLXDhsSOMWPfgbXw; 
				285:VcDzTcOFndjUjhnRfxTN<=VcDzTcOFndjUjhnRfxTN+CHmFHLXDhsSOMWPfgbXw; 
				286:ScSvdbbLcbwcpTKFudIt<=ScSvdbbLcbwcpTKFudIt+CHmFHLXDhsSOMWPfgbXw; 
				287:ZFOGopcNcymIuYXsiiRw<=ZFOGopcNcymIuYXsiiRw+CHmFHLXDhsSOMWPfgbXw; 
				288:zVAojGgdEwSIpPjTZZId<=zVAojGgdEwSIpPjTZZId+CHmFHLXDhsSOMWPfgbXw; 
				289:qwGWpRzKYsDLRvxcxAAH<=qwGWpRzKYsDLRvxcxAAH+CHmFHLXDhsSOMWPfgbXw; 
				290:WPkpODdzyINGGhuwZyoF<=WPkpODdzyINGGhuwZyoF+CHmFHLXDhsSOMWPfgbXw; 
				291:BaxiLnGgFxSKHVKkEWrL<=BaxiLnGgFxSKHVKkEWrL+CHmFHLXDhsSOMWPfgbXw; 
				292:cChsgcLGnvNEmegZREam<=cChsgcLGnvNEmegZREam+CHmFHLXDhsSOMWPfgbXw; 
				293:FRCWHcmIuMUUWgdYMzWu<=FRCWHcmIuMUUWgdYMzWu+CHmFHLXDhsSOMWPfgbXw; 
				294:QDYrIGBlnoXdNCUflHOP<=QDYrIGBlnoXdNCUflHOP+CHmFHLXDhsSOMWPfgbXw; 
				295:zzYTnLgksIjwqZSweXMf<=zzYTnLgksIjwqZSweXMf+CHmFHLXDhsSOMWPfgbXw; 
				296:cWljGAlocPwsnrDyMjHO<=cWljGAlocPwsnrDyMjHO+CHmFHLXDhsSOMWPfgbXw; 
				297:JPYOnWGSGjFuHZfQBaEZ<=JPYOnWGSGjFuHZfQBaEZ+CHmFHLXDhsSOMWPfgbXw; 
				298:VzfYJEwelHYPMpUSDmsC<=VzfYJEwelHYPMpUSDmsC+CHmFHLXDhsSOMWPfgbXw; 
				299:XYQGKDohhXYVCeaCtmre<=XYQGKDohhXYVCeaCtmre+CHmFHLXDhsSOMWPfgbXw; 
				300:GbajCDnxXLGTStnsYsds<=GbajCDnxXLGTStnsYsds+CHmFHLXDhsSOMWPfgbXw; 
				301:THlQvXwjkuLqdcMtPxBy<=THlQvXwjkuLqdcMtPxBy+CHmFHLXDhsSOMWPfgbXw; 
				302:avkJIgYNFpvoyRkxaMTC<=avkJIgYNFpvoyRkxaMTC+CHmFHLXDhsSOMWPfgbXw; 
				303:yhgnNUWIhVDlrtUDGEZn<=yhgnNUWIhVDlrtUDGEZn+CHmFHLXDhsSOMWPfgbXw; 
				304:lHvULbFfwhQgtqfjhwzH<=lHvULbFfwhQgtqfjhwzH+CHmFHLXDhsSOMWPfgbXw; 
				305:TymwlUFeZUaLhFoWTZzU<=TymwlUFeZUaLhFoWTZzU+CHmFHLXDhsSOMWPfgbXw; 
				306:obAWtmAwdFBYPXQlSuSy<=obAWtmAwdFBYPXQlSuSy+CHmFHLXDhsSOMWPfgbXw; 
				307:VBJGcheVZYcxGpvcuBoi<=VBJGcheVZYcxGpvcuBoi+CHmFHLXDhsSOMWPfgbXw; 
				308:NpcOSbiIpOcdgCjboENs<=NpcOSbiIpOcdgCjboENs+CHmFHLXDhsSOMWPfgbXw; 
				309:PiHYPPmDrZQNPnlqBFSt<=PiHYPPmDrZQNPnlqBFSt+CHmFHLXDhsSOMWPfgbXw; 
				310:rOXoAhCRFHntxISYSkye<=rOXoAhCRFHntxISYSkye+CHmFHLXDhsSOMWPfgbXw; 
				311:IsXHeZVJKogNnFFfJwvx<=IsXHeZVJKogNnFFfJwvx+CHmFHLXDhsSOMWPfgbXw; 
				312:BtfuDWbiQheMoNKySKtm<=BtfuDWbiQheMoNKySKtm+CHmFHLXDhsSOMWPfgbXw; 
				313:lsMUeaCgYLjCPUiUXaIc<=lsMUeaCgYLjCPUiUXaIc+CHmFHLXDhsSOMWPfgbXw; 
				314:kTdnGvNmLrhbepFdhZCh<=kTdnGvNmLrhbepFdhZCh+CHmFHLXDhsSOMWPfgbXw; 
				315:vKbnovNlLRioZoJsQunL<=vKbnovNlLRioZoJsQunL+CHmFHLXDhsSOMWPfgbXw; 
				316:nXBrtwwgIArkXUbHKAye<=nXBrtwwgIArkXUbHKAye+CHmFHLXDhsSOMWPfgbXw; 
				317:czvIYhYPaYPpRHUBJMFc<=czvIYhYPaYPpRHUBJMFc+CHmFHLXDhsSOMWPfgbXw; 
				318:nsezjQWxmqwzmxCwosDv<=nsezjQWxmqwzmxCwosDv+CHmFHLXDhsSOMWPfgbXw; 
				319:ruIyZIesSthmxIaXEtrJ<=ruIyZIesSthmxIaXEtrJ+CHmFHLXDhsSOMWPfgbXw; 
				320:cXQjLxPFTWRBhlJmdxUJ<=cXQjLxPFTWRBhlJmdxUJ+CHmFHLXDhsSOMWPfgbXw; 
				321:GPoMmfciZsakCXuJMdbD<=GPoMmfciZsakCXuJMdbD+CHmFHLXDhsSOMWPfgbXw; 
				322:sZUCFycPxeatsZozmHJN<=sZUCFycPxeatsZozmHJN+CHmFHLXDhsSOMWPfgbXw; 
				323:XbnmwpButuNSkogDlbQb<=XbnmwpButuNSkogDlbQb+CHmFHLXDhsSOMWPfgbXw; 
				324:wdkDXnIkWnpQMmswGQeU<=wdkDXnIkWnpQMmswGQeU+CHmFHLXDhsSOMWPfgbXw; 
				325:KpEHEcApUpQBvCLoAeYT<=KpEHEcApUpQBvCLoAeYT+CHmFHLXDhsSOMWPfgbXw; 
				326:KsaghLmgaRvpRfCktbJZ<=KsaghLmgaRvpRfCktbJZ+CHmFHLXDhsSOMWPfgbXw; 
				327:lZVGNfUlVmsuLbJxnQDA<=lZVGNfUlVmsuLbJxnQDA+CHmFHLXDhsSOMWPfgbXw; 
				328:rMBkqrLcKhflEMUYxGkE<=rMBkqrLcKhflEMUYxGkE+CHmFHLXDhsSOMWPfgbXw; 
				329:wMlYFxkSbZTCTvhQOIei<=wMlYFxkSbZTCTvhQOIei+CHmFHLXDhsSOMWPfgbXw; 
				330:WQGVbnQQZGQWVmpcxvbb<=WQGVbnQQZGQWVmpcxvbb+CHmFHLXDhsSOMWPfgbXw; 
				331:AzsKalhmBYUitbArLbcU<=AzsKalhmBYUitbArLbcU+CHmFHLXDhsSOMWPfgbXw; 
				332:ekrMWzROxYoWtRpdbLZH<=ekrMWzROxYoWtRpdbLZH+CHmFHLXDhsSOMWPfgbXw; 
				333:uLMmObkZiwzDlReqMwJN<=uLMmObkZiwzDlReqMwJN+CHmFHLXDhsSOMWPfgbXw; 
				334:eAEEsZkRTlfXOeEdICRO<=eAEEsZkRTlfXOeEdICRO+CHmFHLXDhsSOMWPfgbXw; 
				335:DyXCiZssIzbywKGAbIwY<=DyXCiZssIzbywKGAbIwY+CHmFHLXDhsSOMWPfgbXw; 
				336:wBOVUPcFUWzhOUKDlJVa<=wBOVUPcFUWzhOUKDlJVa+CHmFHLXDhsSOMWPfgbXw; 
				337:BCsgCSHvysHWLteqbRMX<=BCsgCSHvysHWLteqbRMX+CHmFHLXDhsSOMWPfgbXw; 
				338:FrvVghZEElOfAJGPEURk<=FrvVghZEElOfAJGPEURk+CHmFHLXDhsSOMWPfgbXw; 
				339:DHNpdfPdlvcIeMhPYCBD<=DHNpdfPdlvcIeMhPYCBD+CHmFHLXDhsSOMWPfgbXw; 
				340:ByKBiFClfZeeoBwNqVdH<=ByKBiFClfZeeoBwNqVdH+CHmFHLXDhsSOMWPfgbXw; 
				341:muXlkjUrAqYazTUUGcVg<=muXlkjUrAqYazTUUGcVg+CHmFHLXDhsSOMWPfgbXw; 
				342:rZlIolWetZZffpSrlMAn<=rZlIolWetZZffpSrlMAn+CHmFHLXDhsSOMWPfgbXw; 
				343:fCxfzzVrwjVhwiuAOpOD<=fCxfzzVrwjVhwiuAOpOD+CHmFHLXDhsSOMWPfgbXw; 
				344:VHDrEEGVFWccsKXzbEjD<=VHDrEEGVFWccsKXzbEjD+CHmFHLXDhsSOMWPfgbXw; 
				345:pgbmZFwAnGMkExuHZexG<=pgbmZFwAnGMkExuHZexG+CHmFHLXDhsSOMWPfgbXw; 
				346:CYTIFZXRYHDOwAOpYhTY<=CYTIFZXRYHDOwAOpYhTY+CHmFHLXDhsSOMWPfgbXw; 
				347:hzujftnKaamrwjRBenpS<=hzujftnKaamrwjRBenpS+CHmFHLXDhsSOMWPfgbXw; 
				348:DwBiXGPwomcqrFUiwGKO<=DwBiXGPwomcqrFUiwGKO+CHmFHLXDhsSOMWPfgbXw; 
				349:TxOTbaXnfvTWWAEMVKsT<=TxOTbaXnfvTWWAEMVKsT+CHmFHLXDhsSOMWPfgbXw; 
				350:VBPMSBgUzhZWqifRFXLt<=VBPMSBgUzhZWqifRFXLt+CHmFHLXDhsSOMWPfgbXw; 
				351:fBEMznDkaUpJbucpUFUs<=fBEMznDkaUpJbucpUFUs+CHmFHLXDhsSOMWPfgbXw; 
				352:RXuUWWKfwotmzMaIdOHs<=RXuUWWKfwotmzMaIdOHs+CHmFHLXDhsSOMWPfgbXw; 
				353:DScSrBltRCaJuMKRHxjp<=DScSrBltRCaJuMKRHxjp+CHmFHLXDhsSOMWPfgbXw; 
				354:yKhNJjIQvjuuxuKGtNvD<=yKhNJjIQvjuuxuKGtNvD+CHmFHLXDhsSOMWPfgbXw; 
				355:MBLbhXLxXGZHZERKIoYb<=MBLbhXLxXGZHZERKIoYb+CHmFHLXDhsSOMWPfgbXw; 
				356:AiFthZhNPfZiXSnyPCOt<=AiFthZhNPfZiXSnyPCOt+CHmFHLXDhsSOMWPfgbXw; 
				357:uDpYTElkHJsWMgegRIkv<=uDpYTElkHJsWMgegRIkv+CHmFHLXDhsSOMWPfgbXw; 
				358:LqJHECWMJlDdyFDTTZZH<=LqJHECWMJlDdyFDTTZZH+CHmFHLXDhsSOMWPfgbXw; 
				359:ohfsyAOCKLVNdUfnlZGT<=ohfsyAOCKLVNdUfnlZGT+CHmFHLXDhsSOMWPfgbXw; 
				360:MOoDdDePAGBzQbLCZlwX<=MOoDdDePAGBzQbLCZlwX+CHmFHLXDhsSOMWPfgbXw; 
				361:MHLazVdHgoSmGTltAxsJ<=MHLazVdHgoSmGTltAxsJ+CHmFHLXDhsSOMWPfgbXw; 
				362:CYSqcBzpHDXSSATrgQjL<=CYSqcBzpHDXSSATrgQjL+CHmFHLXDhsSOMWPfgbXw; 
				363:rPKZMoWgFDpDSJXXQmEU<=rPKZMoWgFDpDSJXXQmEU+CHmFHLXDhsSOMWPfgbXw; 
				364:hniufLGfdzmHbDIvsTIo<=hniufLGfdzmHbDIvsTIo+CHmFHLXDhsSOMWPfgbXw; 
				365:wTfPVycgpDcgGCOQhJjH<=wTfPVycgpDcgGCOQhJjH+CHmFHLXDhsSOMWPfgbXw; 
				366:lcOMvsbHZmIJccXoDkqZ<=lcOMvsbHZmIJccXoDkqZ+CHmFHLXDhsSOMWPfgbXw; 
				367:UKirjTCurmcGUGGogrnh<=UKirjTCurmcGUGGogrnh+CHmFHLXDhsSOMWPfgbXw; 
				368:KVLRCNcgwgdezgxdbtiz<=KVLRCNcgwgdezgxdbtiz+CHmFHLXDhsSOMWPfgbXw; 
				369:ISUkQBFCDDhkmXDnEdVT<=ISUkQBFCDDhkmXDnEdVT+CHmFHLXDhsSOMWPfgbXw; 
				370:wLiUXxuAUdxCuAoAbUxH<=wLiUXxuAUdxCuAoAbUxH+CHmFHLXDhsSOMWPfgbXw; 
				371:vQNMUmgdbJJDFKzsjqLK<=vQNMUmgdbJJDFKzsjqLK+CHmFHLXDhsSOMWPfgbXw; 
				372:PPaVHoPQXNFqYDIgCroQ<=PPaVHoPQXNFqYDIgCroQ+CHmFHLXDhsSOMWPfgbXw; 
				373:fZmgOJpwMcdeRjEcecxZ<=fZmgOJpwMcdeRjEcecxZ+CHmFHLXDhsSOMWPfgbXw; 
				374:pXxRQDEgUJLwgwAsNvmV<=pXxRQDEgUJLwgwAsNvmV+CHmFHLXDhsSOMWPfgbXw; 
				375:JWyFVCrskBwarfgMzbIK<=JWyFVCrskBwarfgMzbIK+CHmFHLXDhsSOMWPfgbXw; 
				376:nLMIykvKsueQiebJRjaB<=nLMIykvKsueQiebJRjaB+CHmFHLXDhsSOMWPfgbXw; 
				377:MwUAnLVNdEpwKFXarSrE<=MwUAnLVNdEpwKFXarSrE+CHmFHLXDhsSOMWPfgbXw; 
				378:rwKFeNNlWzDutFvKudZd<=rwKFeNNlWzDutFvKudZd+CHmFHLXDhsSOMWPfgbXw; 
				379:YFTuhpacOohGrtlEUgyn<=YFTuhpacOohGrtlEUgyn+CHmFHLXDhsSOMWPfgbXw; 
				380:orsjfJIPQQvjIhvrnfZT<=orsjfJIPQQvjIhvrnfZT+CHmFHLXDhsSOMWPfgbXw; 
				381:beooHOrejCcWcSXDuAMs<=beooHOrejCcWcSXDuAMs+CHmFHLXDhsSOMWPfgbXw; 
				382:wLFqLqnhtGKyjhXVaXLu<=wLFqLqnhtGKyjhXVaXLu+CHmFHLXDhsSOMWPfgbXw; 
				383:VhlEwlgxfirfMpIAJZhE<=VhlEwlgxfirfMpIAJZhE+CHmFHLXDhsSOMWPfgbXw; 
				384:ybSCwixJTEhXYyRpEeDj<=ybSCwixJTEhXYyRpEeDj+CHmFHLXDhsSOMWPfgbXw; 
				385:PLAwknGzfcioZVaFOQCX<=PLAwknGzfcioZVaFOQCX+CHmFHLXDhsSOMWPfgbXw; 
				386:WdDdHRBJZdBPCxmYbWdk<=WdDdHRBJZdBPCxmYbWdk+CHmFHLXDhsSOMWPfgbXw; 
				387:BIxIzsQvWljjGYxMCQtS<=BIxIzsQvWljjGYxMCQtS+CHmFHLXDhsSOMWPfgbXw; 
				388:TZYUrtPvAdyOAezlYVJO<=TZYUrtPvAdyOAezlYVJO+CHmFHLXDhsSOMWPfgbXw; 
				389:qPqZhRZBobhmAXNGrsmh<=qPqZhRZBobhmAXNGrsmh+CHmFHLXDhsSOMWPfgbXw; 
				390:BCGaGkllXBcyohBosHqS<=BCGaGkllXBcyohBosHqS+CHmFHLXDhsSOMWPfgbXw; 
				391:pcgiabuotmBHXKOYDDAq<=pcgiabuotmBHXKOYDDAq+CHmFHLXDhsSOMWPfgbXw; 
				392:VidvAsXIfsppEpKtZeYc<=VidvAsXIfsppEpKtZeYc+CHmFHLXDhsSOMWPfgbXw; 
				393:lGfaCxQtDihDBzWEuyaH<=lGfaCxQtDihDBzWEuyaH+CHmFHLXDhsSOMWPfgbXw; 
				394:ucwrtDfHQDZIjkmTmCvN<=ucwrtDfHQDZIjkmTmCvN+CHmFHLXDhsSOMWPfgbXw; 
				395:dayIzRpYaQRnEjXynbCm<=dayIzRpYaQRnEjXynbCm+CHmFHLXDhsSOMWPfgbXw; 
				396:vqgpItmCwuhiwKZyFXMt<=vqgpItmCwuhiwKZyFXMt+CHmFHLXDhsSOMWPfgbXw; 
				397:FnVEwsGKlXZfUqxZGqHn<=FnVEwsGKlXZfUqxZGqHn+CHmFHLXDhsSOMWPfgbXw; 
				398:bitnzrgsExKEWSXnsRZq<=bitnzrgsExKEWSXnsRZq+CHmFHLXDhsSOMWPfgbXw; 
				399:eYsNwIgUOqnSppAZBKfW<=eYsNwIgUOqnSppAZBKfW+CHmFHLXDhsSOMWPfgbXw; 
				400:FXTNpbkOJRifihZRkFUk<=FXTNpbkOJRifihZRkFUk+CHmFHLXDhsSOMWPfgbXw; 
				401:UCyPKegIVHgIqztViRHP<=UCyPKegIVHgIqztViRHP+CHmFHLXDhsSOMWPfgbXw; 
				402:urwbynurHojveDuzQAqY<=urwbynurHojveDuzQAqY+CHmFHLXDhsSOMWPfgbXw; 
				403:djsdiJHbeUEoOocTIVAL<=djsdiJHbeUEoOocTIVAL+CHmFHLXDhsSOMWPfgbXw; 
				404:juEeWiBDxjlSPOBoDWca<=juEeWiBDxjlSPOBoDWca+CHmFHLXDhsSOMWPfgbXw; 
				405:ZfhQiwfaJoKgwqVVBKhf<=ZfhQiwfaJoKgwqVVBKhf+CHmFHLXDhsSOMWPfgbXw; 
				406:SNnVNrhdPUfxhixiespl<=SNnVNrhdPUfxhixiespl+CHmFHLXDhsSOMWPfgbXw; 
				407:cHHoYqPSIzoxFEuXvNLY<=cHHoYqPSIzoxFEuXvNLY+CHmFHLXDhsSOMWPfgbXw; 
				408:hLpCUWbILJOjqbDhVEwn<=hLpCUWbILJOjqbDhVEwn+CHmFHLXDhsSOMWPfgbXw; 
				409:itXQCyFacJzvPyzfGwVe<=itXQCyFacJzvPyzfGwVe+CHmFHLXDhsSOMWPfgbXw; 
				410:iujmIQQClXPYAKjueUBD<=iujmIQQClXPYAKjueUBD+CHmFHLXDhsSOMWPfgbXw; 
				411:BjdcbpGuKPxnpZzFTfte<=BjdcbpGuKPxnpZzFTfte+CHmFHLXDhsSOMWPfgbXw; 
				412:ZQFzyLJsVraTCGkqQcZA<=ZQFzyLJsVraTCGkqQcZA+CHmFHLXDhsSOMWPfgbXw; 
				413:fADZyEOwTyWvSQFgOnwG<=fADZyEOwTyWvSQFgOnwG+CHmFHLXDhsSOMWPfgbXw; 
				414:xbhqvpXrDTlnyBNQeAlC<=xbhqvpXrDTlnyBNQeAlC+CHmFHLXDhsSOMWPfgbXw; 
				415:usigvHtlPqTHmByMEGLy<=usigvHtlPqTHmByMEGLy+CHmFHLXDhsSOMWPfgbXw; 
				416:EqRnSoIxQaLPlCNmpBmq<=EqRnSoIxQaLPlCNmpBmq+CHmFHLXDhsSOMWPfgbXw; 
				417:VzsEzvUFwafgXDXiMnOI<=VzsEzvUFwafgXDXiMnOI+CHmFHLXDhsSOMWPfgbXw; 
				418:qjQChEpAPSbKmoDGRppN<=qjQChEpAPSbKmoDGRppN+CHmFHLXDhsSOMWPfgbXw; 
				419:XBdmfGxuWrXGMBFOANKF<=XBdmfGxuWrXGMBFOANKF+CHmFHLXDhsSOMWPfgbXw; 
				420:iHWmgCopJntOccGPObxn<=iHWmgCopJntOccGPObxn+CHmFHLXDhsSOMWPfgbXw; 
				421:eeoTbTyuwxPCsjuUGnLj<=eeoTbTyuwxPCsjuUGnLj+CHmFHLXDhsSOMWPfgbXw; 
				422:MkxrURKJtUzHVTfBwhoO<=MkxrURKJtUzHVTfBwhoO+CHmFHLXDhsSOMWPfgbXw; 
				423:USFkaPtDBVOjbGpLXKUX<=USFkaPtDBVOjbGpLXKUX+CHmFHLXDhsSOMWPfgbXw; 
				424:xcBSpPXNgyeMCKwBcsxX<=xcBSpPXNgyeMCKwBcsxX+CHmFHLXDhsSOMWPfgbXw; 
				425:APZhwjfiYOuKluWEaTIj<=APZhwjfiYOuKluWEaTIj+CHmFHLXDhsSOMWPfgbXw; 
				426:eiYeGwmYgODBCzcNuNtn<=eiYeGwmYgODBCzcNuNtn+CHmFHLXDhsSOMWPfgbXw; 
				427:rmoQVcRSrSeskIibJzCc<=rmoQVcRSrSeskIibJzCc+CHmFHLXDhsSOMWPfgbXw; 
				428:AzSDmFqniQGEkrUvtcQd<=AzSDmFqniQGEkrUvtcQd+CHmFHLXDhsSOMWPfgbXw; 
				429:BYQMYRDRDKXGHnLYQyKL<=BYQMYRDRDKXGHnLYQyKL+CHmFHLXDhsSOMWPfgbXw; 
				430:iYaojeeenaSObFkfIEyS<=iYaojeeenaSObFkfIEyS+CHmFHLXDhsSOMWPfgbXw; 
				431:OvjWCALXGQonpSVNSUDx<=OvjWCALXGQonpSVNSUDx+CHmFHLXDhsSOMWPfgbXw; 
				432:QNSQONiKmlvpucXZsAKo<=QNSQONiKmlvpucXZsAKo+CHmFHLXDhsSOMWPfgbXw; 
				433:RKLbOFQSgMkwEdftvnBQ<=RKLbOFQSgMkwEdftvnBQ+CHmFHLXDhsSOMWPfgbXw; 
				434:hoPvrLDkwXFTkYESCUcp<=hoPvrLDkwXFTkYESCUcp+CHmFHLXDhsSOMWPfgbXw; 
				435:hShwACbdYktXmGxyazAM<=hShwACbdYktXmGxyazAM+CHmFHLXDhsSOMWPfgbXw; 
				436:puehHutFkvCRvoGqbSYp<=puehHutFkvCRvoGqbSYp+CHmFHLXDhsSOMWPfgbXw; 
				437:CSpvXCVkXjBnWvAFEiDG<=CSpvXCVkXjBnWvAFEiDG+CHmFHLXDhsSOMWPfgbXw; 
				438:GBnbMGmdJLNqPHpTRJqo<=GBnbMGmdJLNqPHpTRJqo+CHmFHLXDhsSOMWPfgbXw; 
				439:PQFlqUWXvhfFTKRniEDA<=PQFlqUWXvhfFTKRniEDA+CHmFHLXDhsSOMWPfgbXw; 
				440:mNQfwTdWpUOnxIhbTYfU<=mNQfwTdWpUOnxIhbTYfU+CHmFHLXDhsSOMWPfgbXw; 
				441:ldQowZgtPeXlzjFcyWQl<=ldQowZgtPeXlzjFcyWQl+CHmFHLXDhsSOMWPfgbXw; 
				442:HYWHYpKWyjTHzWIzGNeE<=HYWHYpKWyjTHzWIzGNeE+CHmFHLXDhsSOMWPfgbXw; 
				443:vsHmuANStIQsYgoNHsHw<=vsHmuANStIQsYgoNHsHw+CHmFHLXDhsSOMWPfgbXw; 
				444:tYWmIUymjXADFjUmKFpP<=tYWmIUymjXADFjUmKFpP+CHmFHLXDhsSOMWPfgbXw; 
				445:OQmggBTvOqhAXBiDJeaP<=OQmggBTvOqhAXBiDJeaP+CHmFHLXDhsSOMWPfgbXw; 
				446:EFcUAERFHbivPwgHAMQa<=EFcUAERFHbivPwgHAMQa+CHmFHLXDhsSOMWPfgbXw; 
				447:jpbydIYGKyCwhjgemImi<=jpbydIYGKyCwhjgemImi+CHmFHLXDhsSOMWPfgbXw; 
				448:OVYjPuZDVHOTTeuFPkrT<=OVYjPuZDVHOTTeuFPkrT+CHmFHLXDhsSOMWPfgbXw; 
				449:DqhwOfIUxBzsVSgEjWzC<=DqhwOfIUxBzsVSgEjWzC+CHmFHLXDhsSOMWPfgbXw; 
				450:plztNCDwyKBliboMvXKs<=plztNCDwyKBliboMvXKs+CHmFHLXDhsSOMWPfgbXw; 
				451:GojVETmCGfWcYwVYimBv<=GojVETmCGfWcYwVYimBv+CHmFHLXDhsSOMWPfgbXw; 
				452:aogDiFiAXQqphSrsQbJV<=aogDiFiAXQqphSrsQbJV+CHmFHLXDhsSOMWPfgbXw; 
				453:rCOKgSoVLfXaUWFdsBnJ<=rCOKgSoVLfXaUWFdsBnJ+CHmFHLXDhsSOMWPfgbXw; 
				454:ZuONZDcmHxALaUULMEAA<=ZuONZDcmHxALaUULMEAA+CHmFHLXDhsSOMWPfgbXw; 
				455:KIjEeYrBOSrzUMqGYBsV<=KIjEeYrBOSrzUMqGYBsV+CHmFHLXDhsSOMWPfgbXw; 
				456:ZBocacKljeyYorCiQgzQ<=ZBocacKljeyYorCiQgzQ+CHmFHLXDhsSOMWPfgbXw; 
				457:mqazMnBgYnlLqLRzaNYx<=mqazMnBgYnlLqLRzaNYx+CHmFHLXDhsSOMWPfgbXw; 
				458:oyfKvpCwkpoCCxTglCJr<=oyfKvpCwkpoCCxTglCJr+CHmFHLXDhsSOMWPfgbXw; 
				459:NGNEGckWnRLaqnjOKOmx<=NGNEGckWnRLaqnjOKOmx+CHmFHLXDhsSOMWPfgbXw; 
				460:cVWqyzzrUUodYFbrorBz<=cVWqyzzrUUodYFbrorBz+CHmFHLXDhsSOMWPfgbXw; 
				461:RjwugczIYXEQzzmUrnYh<=RjwugczIYXEQzzmUrnYh+CHmFHLXDhsSOMWPfgbXw; 
				462:lEqWgKBWIbLvYwrXeDtN<=lEqWgKBWIbLvYwrXeDtN+CHmFHLXDhsSOMWPfgbXw; 
				463:DhnZhzYLzUMXzuxLMdpR<=DhnZhzYLzUMXzuxLMdpR+CHmFHLXDhsSOMWPfgbXw; 
				464:WwogGcAbNuwPRaXHfllR<=WwogGcAbNuwPRaXHfllR+CHmFHLXDhsSOMWPfgbXw; 
				465:fymbKnqnRYaHIRuPXxle<=fymbKnqnRYaHIRuPXxle+CHmFHLXDhsSOMWPfgbXw; 
				466:nJWkhXEkUmrasSyMThpL<=nJWkhXEkUmrasSyMThpL+CHmFHLXDhsSOMWPfgbXw; 
				467:qXNWBYTrrKKKGSroThrT<=qXNWBYTrrKKKGSroThrT+CHmFHLXDhsSOMWPfgbXw; 
				468:OWgmvdYcTEmvwkEuDkJS<=OWgmvdYcTEmvwkEuDkJS+CHmFHLXDhsSOMWPfgbXw; 
				469:urpaOisfjSiDXEZoTBsG<=urpaOisfjSiDXEZoTBsG+CHmFHLXDhsSOMWPfgbXw; 
				470:mveotDylkopgLZJFFBVl<=mveotDylkopgLZJFFBVl+CHmFHLXDhsSOMWPfgbXw; 
				471:CCXECvtOeIBEOFePtIRw<=CCXECvtOeIBEOFePtIRw+CHmFHLXDhsSOMWPfgbXw; 
				472:iYYwLjjGMjLikfxxrxIB<=iYYwLjjGMjLikfxxrxIB+CHmFHLXDhsSOMWPfgbXw; 
				473:BJhcDugYXUoZuTXYBzJg<=BJhcDugYXUoZuTXYBzJg+CHmFHLXDhsSOMWPfgbXw; 
				474:wpEZHrezpouBVvAiIOpn<=wpEZHrezpouBVvAiIOpn+CHmFHLXDhsSOMWPfgbXw; 
				475:omjfRcaEwaSdXWjgQYUv<=omjfRcaEwaSdXWjgQYUv+CHmFHLXDhsSOMWPfgbXw; 
				476:aWXCrpICnOAsyXgkDTDT<=aWXCrpICnOAsyXgkDTDT+CHmFHLXDhsSOMWPfgbXw; 
				477:HjXRkNnhDmrrYeoZLfga<=HjXRkNnhDmrrYeoZLfga+CHmFHLXDhsSOMWPfgbXw; 
				478:zDWiKpAenkhcNZIBSNiT<=zDWiKpAenkhcNZIBSNiT+CHmFHLXDhsSOMWPfgbXw; 
				479:UfyNbuBOwMXEdumKnlqN<=UfyNbuBOwMXEdumKnlqN+CHmFHLXDhsSOMWPfgbXw; 
				480:LYSwVHbgNGVrAkuDLmxY<=LYSwVHbgNGVrAkuDLmxY+CHmFHLXDhsSOMWPfgbXw;//}}}
			endcase
		end
	end
	always@(*)
	begin
		if(eojmGbYrZBcDvhuhplcn)
		begin
			case(XWSDWJpZwWFziLcqAlai)
				0:aSItvOfWsSQOkHOHMzuM=iGrqtIPPBFPUhGunhSdw;
    			1:aSItvOfWsSQOkHOHMzuM=CZceBwenUmhgWecdrVuw;
    			2:aSItvOfWsSQOkHOHMzuM=FODhltaveISdQIJPBJhJ;
				default:aSItvOfWsSQOkHOHMzuM=0;
			endcase
		end
		else
		begin
			case(XWSDWJpZwWFziLcqAlai)
				0:aSItvOfWsSQOkHOHMzuM=mBUfUweOiYOTkxaNfvqZ;
    			1:aSItvOfWsSQOkHOHMzuM=XCEBnusbPkduEdkiHxFK;
    			2:aSItvOfWsSQOkHOHMzuM=UKLUuuVquDsMMMMhkoJV;
				default:aSItvOfWsSQOkHOHMzuM=0;
			endcase
		end
	end
	always@(*)
	begin
		if(eojmGbYrZBcDvhuhplcn) 
		begin
			case(XWSDWJpZwWFziLcqAlai) 
   				0:kAXRTBBnwMdFccjIlXSw=qUkWgSUxlHDGwaShnpJD;
    			1:kAXRTBBnwMdFccjIlXSw=AKnQHFnRxMsayGvtbpFT;
    			2:kAXRTBBnwMdFccjIlXSw=EdvpzeTpOWEloDTnpLTm;
				default:kAXRTBBnwMdFccjIlXSw=0;
			endcase 
		end
		else
		begin
			case(XWSDWJpZwWFziLcqAlai)
 				0:kAXRTBBnwMdFccjIlXSw=vWFpyuXCRPPETqWnXLgO;
    			1:kAXRTBBnwMdFccjIlXSw=dbsLvjpjMhdBsPiUgbjQ;
    			2:kAXRTBBnwMdFccjIlXSw=oXZLEogkFzslyJXIZmAm;
				default:kAXRTBBnwMdFccjIlXSw=0;
			endcase
		end
	end

	always@(*)
	begin
		if(eojmGbYrZBcDvhuhplcn)
		begin
			case(XWSDWJpZwWFziLcqAlai)
    			0: oEDxWLutHlOkrCgasnsy=RdPhRZcalGKJvMOvrAIh;
    			1: oEDxWLutHlOkrCgasnsy=xMPttPagqqqJUKztQdOZ;
    			2: oEDxWLutHlOkrCgasnsy=YCteCIAKCruidjpeILHG;
  				default:oEDxWLutHlOkrCgasnsy=0;
			endcase
		end
		else
		begin	
			case(XWSDWJpZwWFziLcqAlai)
				0: oEDxWLutHlOkrCgasnsy=nxlEkFPUCwQVbIQJmgbx;
				1: oEDxWLutHlOkrCgasnsy=SVzsQtfHGQqXqNoloxvo;
				2: oEDxWLutHlOkrCgasnsy=vMLEZaXExwsFFvafFmfc;
  				default:oEDxWLutHlOkrCgasnsy=0;
			endcase
		end
	end


	always@(*)
	begin
		if(eojmGbYrZBcDvhuhplcn)
		begin
			case(XWSDWJpZwWFziLcqAlai)
   				0:CHmFHLXDhsSOMWPfgbXw=LkKGICfCcYyYLBJKtucQ;
    			1:CHmFHLXDhsSOMWPfgbXw=SupobFuabxSWuLFQTEEe;
    			2:CHmFHLXDhsSOMWPfgbXw=BUOYkUPXSUGjGnnMOiLz;
				default:CHmFHLXDhsSOMWPfgbXw=0;
			endcase
		end
		else
		begin
			case(XWSDWJpZwWFziLcqAlai)
 				0:CHmFHLXDhsSOMWPfgbXw=tOmHmkYobOhcasHrvveC;
    			1:CHmFHLXDhsSOMWPfgbXw=HMRNTVVBwfsQwiaIOdeu;
    			2:CHmFHLXDhsSOMWPfgbXw=hGCZylpOryFfZNhxLZOH;
				default:CHmFHLXDhsSOMWPfgbXw=0;
			endcase
		end
	end

	always@(posedge rd_clk or negedge rst)
	begin
	    if(!rst)
			bVNTszDvPimBrKwNycBW<=0;
		else if(rst_syn)
			bVNTszDvPimBrKwNycBW<=0;
		else if(gStNdqadtalDMswfRuqW==CAL_SLOPE_1)     
		begin
			if(TLXWChymSkORZZFunpRb)
				bVNTszDvPimBrKwNycBW<=480;
			else
				bVNTszDvPimBrKwNycBW<=qaVKoOckmCbhBtxSbviM+(ARQLJGuTZBnFJHXDoAkT<<4);
		end
	end
	always@(posedge rd_clk or negedge rst)
	begin
	    if(!rst) 
			CTJvELJpTGwHTCgirGVs<=0;
		else if(rst_syn)
			CTJvELJpTGwHTCgirGVs<=0;
		else if(gStNdqadtalDMswfRuqW==CAL_SLOPE_2)            
		begin
			if(TLXWChymSkORZZFunpRb)
				CTJvELJpTGwHTCgirGVs<=0;
			else CTJvELJpTGwHTCgirGVs<=qaVKoOckmCbhBtxSbviM+(ARQLJGuTZBnFJHXDoAkT<<4);
		end
	end
	always@(posedge rd_clk or negedge rst)
	begin
	    if(!rst)
			OhIQvlSNredlAvEzVwlD<=0;
		else if(rst_syn)
			OhIQvlSNredlAvEzVwlD<=0;
		else if(gStNdqadtalDMswfRuqW==PASS_OVER)
			OhIQvlSNredlAvEzVwlD<=0;
		else if(gStNdqadtalDMswfRuqW==CAL_SLOPE_3)
		begin
			if(bVNTszDvPimBrKwNycBW>=CTJvELJpTGwHTCgirGVs)      
				OhIQvlSNredlAvEzVwlD<=bVNTszDvPimBrKwNycBW-CTJvELJpTGwHTCgirGVs;
			else OhIQvlSNredlAvEzVwlD<=0;                               //
		end
	end


	
	always@(posedge wr_clk or negedge rst)
	begin
	    if(!rst) 
		begin
			RdPhRZcalGKJvMOvrAIh<=0;  
			xMPttPagqqqJUKztQdOZ<=0;
			YCteCIAKCruidjpeILHG<=0;
			nxlEkFPUCwQVbIQJmgbx<=0;
			SVzsQtfHGQqXqNoloxvo<=0;
			vMLEZaXExwsFFvafFmfc<=0;
		end
		else if(rst_syn)
		begin			
			RdPhRZcalGKJvMOvrAIh<=0;  
			xMPttPagqqqJUKztQdOZ<=0;
			YCteCIAKCruidjpeILHG<=0;
			nxlEkFPUCwQVbIQJmgbx<=0;
			SVzsQtfHGQqXqNoloxvo<=0;
			vMLEZaXExwsFFvafFmfc<=0;
		end
		else if(flush_over)
		begin
			if(!eojmGbYrZBcDvhuhplcn)
			begin
				RdPhRZcalGKJvMOvrAIh<=pass_error_plane_sp;
				xMPttPagqqqJUKztQdOZ<=pass_error_plane_mp;
				YCteCIAKCruidjpeILHG<=pass_error_plane_cp;
			end
			else 
			begin
				nxlEkFPUCwQVbIQJmgbx<=pass_error_plane_sp;
				SVzsQtfHGQqXqNoloxvo<=pass_error_plane_mp;
				vMLEZaXExwsFFvafFmfc<=pass_error_plane_cp;
			end
		end



	end
	
	always@(*)
	begin
	    case(wKozjyqvbxpraCSNGCJY)
			0  :  qaVKoOckmCbhBtxSbviM=0 ; //{{{
			1  :  qaVKoOckmCbhBtxSbviM=0 ;
			2  :  qaVKoOckmCbhBtxSbviM=0 ;
			3  :  qaVKoOckmCbhBtxSbviM=0 ;
			4  :  qaVKoOckmCbhBtxSbviM=0 ;
			5  :  qaVKoOckmCbhBtxSbviM=0 ;
			6  :  qaVKoOckmCbhBtxSbviM=1 ;
			7  :  qaVKoOckmCbhBtxSbviM=1 ;
			8  :  qaVKoOckmCbhBtxSbviM=1 ;
			9  :  qaVKoOckmCbhBtxSbviM=1 ;
			10 :  qaVKoOckmCbhBtxSbviM=1 ;
			11 :  qaVKoOckmCbhBtxSbviM=1 ;
			12 :  qaVKoOckmCbhBtxSbviM=1 ;
			13 :  qaVKoOckmCbhBtxSbviM=1 ;
			14 :  qaVKoOckmCbhBtxSbviM=1 ;
			15 :  qaVKoOckmCbhBtxSbviM=1 ;
			16 :  qaVKoOckmCbhBtxSbviM=1 ;
			17 :  qaVKoOckmCbhBtxSbviM=1 ;
			18 :  qaVKoOckmCbhBtxSbviM=2 ;
			19 :  qaVKoOckmCbhBtxSbviM=2 ;
			20 :  qaVKoOckmCbhBtxSbviM=2 ;
			21 :  qaVKoOckmCbhBtxSbviM=2 ;
			22 :  qaVKoOckmCbhBtxSbviM=2 ;
			23 :  qaVKoOckmCbhBtxSbviM=2 ;
			24 :  qaVKoOckmCbhBtxSbviM=2 ;
			25 :  qaVKoOckmCbhBtxSbviM=2 ;
			26 :  qaVKoOckmCbhBtxSbviM=2 ;
			27 :  qaVKoOckmCbhBtxSbviM=2 ;
			28 :  qaVKoOckmCbhBtxSbviM=2 ;
			29 :  qaVKoOckmCbhBtxSbviM=2 ;
			30 :  qaVKoOckmCbhBtxSbviM=3 ;
			31 :  qaVKoOckmCbhBtxSbviM=3 ;
			32 :  qaVKoOckmCbhBtxSbviM=3 ;
			33 :  qaVKoOckmCbhBtxSbviM=3 ;
			34 :  qaVKoOckmCbhBtxSbviM=3 ;
			35 :  qaVKoOckmCbhBtxSbviM=3 ;
			36 :  qaVKoOckmCbhBtxSbviM=3 ;
			37 :  qaVKoOckmCbhBtxSbviM=3 ;
			38 :  qaVKoOckmCbhBtxSbviM=3 ;
			39 :  qaVKoOckmCbhBtxSbviM=3 ;
			40 :  qaVKoOckmCbhBtxSbviM=3 ;
			41 :  qaVKoOckmCbhBtxSbviM=3 ;
			42 :  qaVKoOckmCbhBtxSbviM=4 ;
			43 :  qaVKoOckmCbhBtxSbviM=4 ;
			44 :  qaVKoOckmCbhBtxSbviM=4 ;
			45 :  qaVKoOckmCbhBtxSbviM=4 ;
			46 :  qaVKoOckmCbhBtxSbviM=4 ;
			47 :  qaVKoOckmCbhBtxSbviM=4 ;
			48 :  qaVKoOckmCbhBtxSbviM=4 ;
			49 :  qaVKoOckmCbhBtxSbviM=4 ;
			50 :  qaVKoOckmCbhBtxSbviM=4 ;
			51 :  qaVKoOckmCbhBtxSbviM=4 ;
			52 :  qaVKoOckmCbhBtxSbviM=4 ;
			53 :  qaVKoOckmCbhBtxSbviM=4 ;
			54 :  qaVKoOckmCbhBtxSbviM=4 ;
			55 :  qaVKoOckmCbhBtxSbviM=4 ;
			56 :  qaVKoOckmCbhBtxSbviM=5 ;
			57 :  qaVKoOckmCbhBtxSbviM=5 ;
			58 :  qaVKoOckmCbhBtxSbviM=5 ;
			59 :  qaVKoOckmCbhBtxSbviM=5 ;
			60 :  qaVKoOckmCbhBtxSbviM=5 ;
			61 :  qaVKoOckmCbhBtxSbviM=5 ;
			62 :  qaVKoOckmCbhBtxSbviM=5 ;
			63 :  qaVKoOckmCbhBtxSbviM=5 ;
			64 :  qaVKoOckmCbhBtxSbviM=5 ;
			65 :  qaVKoOckmCbhBtxSbviM=5 ;
			66 :  qaVKoOckmCbhBtxSbviM=5 ;
			67 :  qaVKoOckmCbhBtxSbviM=5 ;
			68 :  qaVKoOckmCbhBtxSbviM=5 ;
			69 :  qaVKoOckmCbhBtxSbviM=6 ;
			70 :  qaVKoOckmCbhBtxSbviM=6 ;
			71 :  qaVKoOckmCbhBtxSbviM=6 ;
			72 :  qaVKoOckmCbhBtxSbviM=6 ;
			73 :  qaVKoOckmCbhBtxSbviM=6 ;
			74 :  qaVKoOckmCbhBtxSbviM=6 ;
			75 :  qaVKoOckmCbhBtxSbviM=6 ;
			76 :  qaVKoOckmCbhBtxSbviM=6 ;
			77 :  qaVKoOckmCbhBtxSbviM=6 ;
			78 :  qaVKoOckmCbhBtxSbviM=6 ;
			79 :  qaVKoOckmCbhBtxSbviM=6 ;
			80 :  qaVKoOckmCbhBtxSbviM=6 ;
			81 :  qaVKoOckmCbhBtxSbviM=6 ;
			82 :  qaVKoOckmCbhBtxSbviM=6 ;
			83 :  qaVKoOckmCbhBtxSbviM=6 ;
			84 :  qaVKoOckmCbhBtxSbviM=7 ;
			85 :  qaVKoOckmCbhBtxSbviM=7 ;
			86 :  qaVKoOckmCbhBtxSbviM=7 ;
			87 :  qaVKoOckmCbhBtxSbviM=7 ;
			88 :  qaVKoOckmCbhBtxSbviM=7 ;
			89 :  qaVKoOckmCbhBtxSbviM=7 ;
			90 :  qaVKoOckmCbhBtxSbviM=7 ;
			91 :  qaVKoOckmCbhBtxSbviM=7 ;
			92 :  qaVKoOckmCbhBtxSbviM=7 ;
			93 :  qaVKoOckmCbhBtxSbviM=7 ;
			94 :  qaVKoOckmCbhBtxSbviM=7 ;
			95 :  qaVKoOckmCbhBtxSbviM=7 ;
			96 :  qaVKoOckmCbhBtxSbviM=7 ;
			97 :  qaVKoOckmCbhBtxSbviM=7 ;
			98 :  qaVKoOckmCbhBtxSbviM=7 ;
			99 :  qaVKoOckmCbhBtxSbviM=8 ;
			100:  qaVKoOckmCbhBtxSbviM=8 ;
			101:  qaVKoOckmCbhBtxSbviM=8 ;
			102:  qaVKoOckmCbhBtxSbviM=8 ;
			103:  qaVKoOckmCbhBtxSbviM=8 ;
			104:  qaVKoOckmCbhBtxSbviM=8 ;
			105:  qaVKoOckmCbhBtxSbviM=8 ;
			106:  qaVKoOckmCbhBtxSbviM=8 ;
			107:  qaVKoOckmCbhBtxSbviM=8 ;
			108:  qaVKoOckmCbhBtxSbviM=8 ;
			109:  qaVKoOckmCbhBtxSbviM=8 ;
			110:  qaVKoOckmCbhBtxSbviM=8 ;
			111:  qaVKoOckmCbhBtxSbviM=8 ;
			112:  qaVKoOckmCbhBtxSbviM=8 ;
			113:  qaVKoOckmCbhBtxSbviM=8 ;
			114:  qaVKoOckmCbhBtxSbviM=9 ;
			115:  qaVKoOckmCbhBtxSbviM=9 ;
			116:  qaVKoOckmCbhBtxSbviM=9 ;
			117:  qaVKoOckmCbhBtxSbviM=9 ;
			118:  qaVKoOckmCbhBtxSbviM=9 ;
			119:  qaVKoOckmCbhBtxSbviM=9 ;
			120:  qaVKoOckmCbhBtxSbviM=9 ;
			121:  qaVKoOckmCbhBtxSbviM=9 ;
			122:  qaVKoOckmCbhBtxSbviM=9 ;
			123:  qaVKoOckmCbhBtxSbviM=9 ;
			124:  qaVKoOckmCbhBtxSbviM=9 ;
			125:  qaVKoOckmCbhBtxSbviM=9 ;
			126:  qaVKoOckmCbhBtxSbviM=9 ;
			127:  qaVKoOckmCbhBtxSbviM=9 ;
			128:  qaVKoOckmCbhBtxSbviM=9 ;  
			129:  qaVKoOckmCbhBtxSbviM=9 ;   
			130:  qaVKoOckmCbhBtxSbviM=9 ;   
			131:  qaVKoOckmCbhBtxSbviM=10;   
			132:  qaVKoOckmCbhBtxSbviM=10;   
			133:  qaVKoOckmCbhBtxSbviM=10;   
			134:  qaVKoOckmCbhBtxSbviM=10;   
			135:  qaVKoOckmCbhBtxSbviM=10;   
			136:  qaVKoOckmCbhBtxSbviM=10;   
			137:  qaVKoOckmCbhBtxSbviM=10;   
			138:  qaVKoOckmCbhBtxSbviM=10;   
			139:  qaVKoOckmCbhBtxSbviM=10;   
			140:  qaVKoOckmCbhBtxSbviM=10;   
			141:  qaVKoOckmCbhBtxSbviM=10;   
			142:  qaVKoOckmCbhBtxSbviM=10;   
			143:  qaVKoOckmCbhBtxSbviM=10;   
			144:  qaVKoOckmCbhBtxSbviM=10;   
			145:  qaVKoOckmCbhBtxSbviM=10;   
			146:  qaVKoOckmCbhBtxSbviM=10;   
			147:  qaVKoOckmCbhBtxSbviM=10;   
			148:  qaVKoOckmCbhBtxSbviM=11;   
			149:  qaVKoOckmCbhBtxSbviM=11;   
			150:  qaVKoOckmCbhBtxSbviM=11;   
			151:  qaVKoOckmCbhBtxSbviM=11;   
			152:  qaVKoOckmCbhBtxSbviM=11;   
			153:  qaVKoOckmCbhBtxSbviM=11;   
			154:  qaVKoOckmCbhBtxSbviM=11;   
			155:  qaVKoOckmCbhBtxSbviM=11;   
			156:  qaVKoOckmCbhBtxSbviM=11;   
			157:  qaVKoOckmCbhBtxSbviM=11;   
			158:  qaVKoOckmCbhBtxSbviM=11;   
			159:  qaVKoOckmCbhBtxSbviM=11;   
			160:  qaVKoOckmCbhBtxSbviM=11;   
			161:  qaVKoOckmCbhBtxSbviM=11;   
			162:  qaVKoOckmCbhBtxSbviM=11;   
			163:  qaVKoOckmCbhBtxSbviM=11;   
			164:  qaVKoOckmCbhBtxSbviM=11;   
			165:  qaVKoOckmCbhBtxSbviM=11;   
			166:  qaVKoOckmCbhBtxSbviM=12;   
			167:  qaVKoOckmCbhBtxSbviM=12;   
			168:  qaVKoOckmCbhBtxSbviM=12;   
			169:  qaVKoOckmCbhBtxSbviM=12;   
			170:  qaVKoOckmCbhBtxSbviM=12;   
			171:  qaVKoOckmCbhBtxSbviM=12;   
			172:  qaVKoOckmCbhBtxSbviM=12;   
			173:  qaVKoOckmCbhBtxSbviM=12;   
			174:  qaVKoOckmCbhBtxSbviM=12;   
			175:  qaVKoOckmCbhBtxSbviM=12;   
			176:  qaVKoOckmCbhBtxSbviM=12;   
			177:  qaVKoOckmCbhBtxSbviM=12;   
			178:  qaVKoOckmCbhBtxSbviM=12;   
			179:  qaVKoOckmCbhBtxSbviM=12;   
			180:  qaVKoOckmCbhBtxSbviM=12;   
			181:  qaVKoOckmCbhBtxSbviM=12;   
			182:  qaVKoOckmCbhBtxSbviM=12;   
			183:  qaVKoOckmCbhBtxSbviM=12;   
			184:  qaVKoOckmCbhBtxSbviM=13;   
			185:  qaVKoOckmCbhBtxSbviM=13;   
			186:  qaVKoOckmCbhBtxSbviM=13;   
			187:  qaVKoOckmCbhBtxSbviM=13;   
			188:  qaVKoOckmCbhBtxSbviM=13;   
			189:  qaVKoOckmCbhBtxSbviM=13;   
			190:  qaVKoOckmCbhBtxSbviM=13;   
			191:  qaVKoOckmCbhBtxSbviM=13;   
			192:  qaVKoOckmCbhBtxSbviM=13;   
			193:  qaVKoOckmCbhBtxSbviM=13;   
			194:  qaVKoOckmCbhBtxSbviM=13;   
			195:  qaVKoOckmCbhBtxSbviM=13;   
			196:  qaVKoOckmCbhBtxSbviM=13;   
			197:  qaVKoOckmCbhBtxSbviM=13;   
			198:  qaVKoOckmCbhBtxSbviM=13;   
			199:  qaVKoOckmCbhBtxSbviM=13;   
			200:  qaVKoOckmCbhBtxSbviM=13;   
			201:  qaVKoOckmCbhBtxSbviM=13;   
			202:  qaVKoOckmCbhBtxSbviM=13;   
			203:  qaVKoOckmCbhBtxSbviM=13;   
			204:  qaVKoOckmCbhBtxSbviM=14;   
			205:  qaVKoOckmCbhBtxSbviM=14;   
			206:  qaVKoOckmCbhBtxSbviM=14;   
			207:  qaVKoOckmCbhBtxSbviM=14;   
			208:  qaVKoOckmCbhBtxSbviM=14;   
			209:  qaVKoOckmCbhBtxSbviM=14;   
			210:  qaVKoOckmCbhBtxSbviM=14;   
			211:  qaVKoOckmCbhBtxSbviM=14;   
			212:  qaVKoOckmCbhBtxSbviM=14;   
			213:  qaVKoOckmCbhBtxSbviM=14;   
			214:  qaVKoOckmCbhBtxSbviM=14;   
			215:  qaVKoOckmCbhBtxSbviM=14;   
			216:  qaVKoOckmCbhBtxSbviM=14;   
			217:  qaVKoOckmCbhBtxSbviM=14;   
			218:  qaVKoOckmCbhBtxSbviM=14;   
			219:  qaVKoOckmCbhBtxSbviM=14;   
			220:  qaVKoOckmCbhBtxSbviM=14;   
			221:  qaVKoOckmCbhBtxSbviM=14;   
			222:  qaVKoOckmCbhBtxSbviM=14;   
			223:  qaVKoOckmCbhBtxSbviM=14;   
			224:  qaVKoOckmCbhBtxSbviM=15;   
			225:  qaVKoOckmCbhBtxSbviM=15;   
			226:  qaVKoOckmCbhBtxSbviM=15;   
			227:  qaVKoOckmCbhBtxSbviM=15;   
			228:  qaVKoOckmCbhBtxSbviM=15;   
			229:  qaVKoOckmCbhBtxSbviM=15;   
			230:  qaVKoOckmCbhBtxSbviM=15;   
			231:  qaVKoOckmCbhBtxSbviM=15;   
			232:  qaVKoOckmCbhBtxSbviM=15;   
			233:  qaVKoOckmCbhBtxSbviM=15;   
			234:  qaVKoOckmCbhBtxSbviM=15;   
			235:  qaVKoOckmCbhBtxSbviM=15;   
			236:  qaVKoOckmCbhBtxSbviM=15;   
			237:  qaVKoOckmCbhBtxSbviM=15;   
			238:  qaVKoOckmCbhBtxSbviM=15;   
			239:  qaVKoOckmCbhBtxSbviM=15;   
			240:  qaVKoOckmCbhBtxSbviM=15;   
			241:  qaVKoOckmCbhBtxSbviM=15;   
			242:  qaVKoOckmCbhBtxSbviM=15;   
			243:  qaVKoOckmCbhBtxSbviM=15;   
			244:  qaVKoOckmCbhBtxSbviM=15;   
			245:  qaVKoOckmCbhBtxSbviM=15;   
			246:  qaVKoOckmCbhBtxSbviM=16;   
			247:  qaVKoOckmCbhBtxSbviM=16;   
			248:  qaVKoOckmCbhBtxSbviM=16;   
			249:  qaVKoOckmCbhBtxSbviM=16;   
			250:  qaVKoOckmCbhBtxSbviM=16;   
			251:  qaVKoOckmCbhBtxSbviM=16;   
			252:  qaVKoOckmCbhBtxSbviM=16;   
			253:  qaVKoOckmCbhBtxSbviM=16;   
			254:  qaVKoOckmCbhBtxSbviM=16;   
			255:  qaVKoOckmCbhBtxSbviM=16;   //}}}
			default:qaVKoOckmCbhBtxSbviM=0 ;
		endcase
	end

	always@(*)
	begin
	    case(gStNdqadtalDMswfRuqW)
			CAL_SLOPE_1:wKozjyqvbxpraCSNGCJY=FssIYlUsXIkosBplffKR;
			CAL_SLOPE_2:wKozjyqvbxpraCSNGCJY=fvbJniljSNczcXeDYDTv;
			default:wKozjyqvbxpraCSNGCJY=0;
		endcase
	end

	always@(posedge rd_clk or negedge rst)
	begin
	    if(!rst)
			XWSDWJpZwWFziLcqAlai<=0;
		else if(rst_syn)
			XWSDWJpZwWFziLcqAlai<=0;
		else 
			begin
				case(gStNdqadtalDMswfRuqW)
					FIND_FIRST_PASS:
					begin
						case(irdAYQxVjzyKmWopQQGP)
							3'b111:XWSDWJpZwWFziLcqAlai<=3;
							3'b110:XWSDWJpZwWFziLcqAlai<=2;
							3'b100:XWSDWJpZwWFziLcqAlai<=1;
							3'b000:XWSDWJpZwWFziLcqAlai<=0;
						endcase                                                     
					end
					NEXT_PASS:XWSDWJpZwWFziLcqAlai<=XWSDWJpZwWFziLcqAlai+1;
					PASS_OVER:XWSDWJpZwWFziLcqAlai<=0;
				endcase
			end

	end

	always@(posedge wr_clk or negedge rst)
	begin
	    if(!rst) 
			eojmGbYrZBcDvhuhplcn<=0;
		else if(rst_syn)
			eojmGbYrZBcDvhuhplcn<=0;
		else if(flush_over)
			eojmGbYrZBcDvhuhplcn<=!eojmGbYrZBcDvhuhplcn;
	end
	
	assign TLXWChymSkORZZFunpRb=(oEDxWLutHlOkrCgasnsy==0)&&(XWSDWJpZwWFziLcqAlai!=3);
	assign FuMFDshlwPAZNriIzdKA=codeblock_counter==15;  
	assign ytSqxoZpMDkNRuAUbZDc=GVfnzKKftzXfxeBqPQMD>=target_byte_number;
	assign nhadPSkgCafxNJCdwkKp=LrLbKGgLtBSEzbICsDNb?2'b10:2'b01;
	assign jMCVmjFKEszeMFGJPhDT=(gStNdqadtalDMswfRuqW==CAL_TRUNCATION_POINT)&&(!ytSqxoZpMDkNRuAUbZDc);
	wire [4:0]yolIhRYCHLHAYQZvudWh=(30-ARQLJGuTZBnFJHXDoAkT);
	assign CxvpyAhqMqQXTLpXgdOB=OHenhlDjGfxNrcoKTDTe<<yolIhRYCHLHAYQZvudWh;
	assign JBFuaKfGSzMztOCsXGjt=rczbRGCFDOHKNTiwObwc<<yolIhRYCHLHAYQZvudWh;
	assign fvbJniljSNczcXeDYDTv=CxvpyAhqMqQXTLpXgdOB[37:30];
	assign FssIYlUsXIkosBplffKR=JBFuaKfGSzMztOCsXGjt[37:30];
	assign OHenhlDjGfxNrcoKTDTe={22'b0,CHmFHLXDhsSOMWPfgbXw[7:0],8'b0};
	assign rczbRGCFDOHKNTiwObwc={oEDxWLutHlOkrCgasnsy,8'b0};
	assign uoqQSqkDyZwtvuETruXA={qUkWgSUxlHDGwaShnpJD,AKnQHFnRxMsayGvtbpFT,EdvpzeTpOWEloDTnpLTm};
	assign AnaDOfYtVBlpyqvNRuwL={vWFpyuXCRPPETqWnXLgO,dbsLvjpjMhdBsPiUgbjQ,oXZLEogkFzslyJXIZmAm};
	assign irdAYQxVjzyKmWopQQGP=eojmGbYrZBcDvhuhplcn?uoqQSqkDyZwtvuETruXA:AnaDOfYtVBlpyqvNRuwL;
	assign GVEVAzxUWjnkLWGcHbCC=(XWSDWJpZwWFziLcqAlai==0)&&(gStNdqadtalDMswfRuqW==SHIFT_PASS_SECOND_HEADER||gStNdqadtalDMswfRuqW==SHIFT_CODESTREAM)&&!qUkWgSUxlHDGwaShnpJD&&eojmGbYrZBcDvhuhplcn;
	assign artgRMUHHAMMXysfVQxf=(XWSDWJpZwWFziLcqAlai==0)&&(gStNdqadtalDMswfRuqW==SHIFT_PASS_SECOND_HEADER||gStNdqadtalDMswfRuqW==SHIFT_CODESTREAM)&&!vWFpyuXCRPPETqWnXLgO&&(!eojmGbYrZBcDvhuhplcn);   
	assign ZOkiujEkXjtpgkcONTax=(XWSDWJpZwWFziLcqAlai==1)&&(gStNdqadtalDMswfRuqW==SHIFT_PASS_SECOND_HEADER||gStNdqadtalDMswfRuqW==SHIFT_CODESTREAM)&&!AKnQHFnRxMsayGvtbpFT&&eojmGbYrZBcDvhuhplcn;
	assign CcBPKbMCVTPpuzcHaNNl=(XWSDWJpZwWFziLcqAlai==1)&&(gStNdqadtalDMswfRuqW==SHIFT_PASS_SECOND_HEADER||gStNdqadtalDMswfRuqW==SHIFT_CODESTREAM)&&!dbsLvjpjMhdBsPiUgbjQ&&(!eojmGbYrZBcDvhuhplcn);   
	assign QcQmUnoklSTURFcjjsxj=(XWSDWJpZwWFziLcqAlai==2)&&(gStNdqadtalDMswfRuqW==SHIFT_PASS_SECOND_HEADER||gStNdqadtalDMswfRuqW==SHIFT_CODESTREAM)&&!EdvpzeTpOWEloDTnpLTm&&eojmGbYrZBcDvhuhplcn;
	assign MQgLtHVUbOxalviVAmNV=(XWSDWJpZwWFziLcqAlai==2)&&(gStNdqadtalDMswfRuqW==SHIFT_PASS_SECOND_HEADER||gStNdqadtalDMswfRuqW==SHIFT_CODESTREAM)&&!oXZLEogkFzslyJXIZmAm&&(!eojmGbYrZBcDvhuhplcn);   


	always@(posedge rd_clk or negedge rst)
	begin
	    if(!rst) 
			gStNdqadtalDMswfRuqW<=tqCfMxDxNMUeAVjaKWqL;
		else if(rst_syn)
			gStNdqadtalDMswfRuqW<=tqCfMxDxNMUeAVjaKWqL;
		else gStNdqadtalDMswfRuqW<=euqWRDzuVBfSvNZlbygs;
	end

	always@(*)
	begin
	    case(gStNdqadtalDMswfRuqW) 
			tqCfMxDxNMUeAVjaKWqL: 
			begin
				if(cal_truncation_point_start) 
					euqWRDzuVBfSvNZlbygs=CAL_TRUNCATION_POINT;
				else if(flush_over)
					euqWRDzuVBfSvNZlbygs=WAITING_WRITE_OVER;	
				else if(one_codeblock_over&&XtrJUtwJnzBPPMzRDosc==0||daVvNjfwJBQRozThYCld!=0 || (nQAnZVgoKyprBQAdRCfA&&(!wEtGDzRjafclnvKxgCSP)))
					euqWRDzuVBfSvNZlbygs=FIND_FIRST_PASS;
				else if(FuMFDshlwPAZNriIzdKA&&codeblock_shift_over)
					euqWRDzuVBfSvNZlbygs=SHIFT_OVER_FLAG;
				else euqWRDzuVBfSvNZlbygs=tqCfMxDxNMUeAVjaKWqL;
			end
			WAITING_WRITE_OVER:
			begin
				if(YfuArrGnpBUyrJxEvVgI==5)
					euqWRDzuVBfSvNZlbygs=FIND_FIRST_PASS;
				else euqWRDzuVBfSvNZlbygs=WAITING_WRITE_OVER;
			end
			FIND_FIRST_PASS:
				begin
					if(XtrJUtwJnzBPPMzRDosc==0||codeblock_shift_over!=0)
						euqWRDzuVBfSvNZlbygs=SHIFT_PASS_FIRST_HEADER;
					else
						euqWRDzuVBfSvNZlbygs=CAL_SLOPE_1;
				end
			CAL_SLOPE_1:euqWRDzuVBfSvNZlbygs=CAL_SLOPE_2;
			CAL_SLOPE_2:euqWRDzuVBfSvNZlbygs=CAL_SLOPE_3;
			CAL_SLOPE_3:euqWRDzuVBfSvNZlbygs=SHIFT_PASS_FIRST_HEADER;
			SHIFT_PASS_FIRST_HEADER:euqWRDzuVBfSvNZlbygs=SHIFT_PASS_SECOND_HEADER;
			SHIFT_PASS_SECOND_HEADER:
				begin
					if(XWSDWJpZwWFziLcqAlai==3)
					begin
						if(daVvNjfwJBQRozThYCld!=0&&(!nQAnZVgoKyprBQAdRCfA))
							euqWRDzuVBfSvNZlbygs=ONE_EMPTY_CODEBLOCK_OVER;
						else
							euqWRDzuVBfSvNZlbygs=PASS_OVER;
					end 
					else euqWRDzuVBfSvNZlbygs=SHIFT_CODESTREAM;
				end
			SHIFT_CODESTREAM:
			begin
				if(kAXRTBBnwMdFccjIlXSw)
				begin
					if(XWSDWJpZwWFziLcqAlai==2||XWSDWJpZwWFziLcqAlai==3)
					begin
						euqWRDzuVBfSvNZlbygs=PASS_OVER;
					end
					else euqWRDzuVBfSvNZlbygs=NEXT_PASS;
				end
				else euqWRDzuVBfSvNZlbygs=SHIFT_CODESTREAM;
			end
			SHIFT_OVER_FLAG:
				euqWRDzuVBfSvNZlbygs=tqCfMxDxNMUeAVjaKWqL;
			NEXT_PASS:euqWRDzuVBfSvNZlbygs=CAL_SLOPE_1;
			PASS_OVER:euqWRDzuVBfSvNZlbygs=tqCfMxDxNMUeAVjaKWqL;
			CAL_TRUNCATION_POINT:
			begin
				if(ytSqxoZpMDkNRuAUbZDc||(jMCVmjFKEszeMFGJPhDT&&lram_address_wr==480))
					euqWRDzuVBfSvNZlbygs=CAL_TRUNCATION_POINT_OVER;
				else euqWRDzuVBfSvNZlbygs=CAL_TRUNCATION_POINT;
			end
			CAL_TRUNCATION_POINT_OVER:euqWRDzuVBfSvNZlbygs=BUFFER;
			BUFFER:euqWRDzuVBfSvNZlbygs=tqCfMxDxNMUeAVjaKWqL;
			ONE_EMPTY_CODEBLOCK_OVER: 
			begin
				if(daVvNjfwJBQRozThYCld==1&&FuMFDshlwPAZNriIzdKA)
					euqWRDzuVBfSvNZlbygs=SHIFT_OVER_FLAG;
				else euqWRDzuVBfSvNZlbygs=tqCfMxDxNMUeAVjaKWqL;
			end 
			default:euqWRDzuVBfSvNZlbygs=tqCfMxDxNMUeAVjaKWqL;
		endcase
	end
	
	fifo_bitplane_256_16	fifo_bitplane (
		.rd_clk			(rd_clk), 
		.wr_clk			(wr_clk),
		.rst_syn			(rst_syn),
		.din			(data_from_mq),
		.pass			(pass_plane),
		.fifo_group		(eojmGbYrZBcDvhuhplcn),
		.rd_data_count_sp_0(LkKGICfCcYyYLBJKtucQ), 
		.rd_data_count_mp_0(SupobFuabxSWuLFQTEEe),
		.rd_data_count_cp_0(BUOYkUPXSUGjGnnMOiLz),
		.rd_data_count_sp_1(tOmHmkYobOhcasHrvveC),
		.rd_data_count_mp_1(HMRNTVVBwfsQwiaIOdeu),
		.rd_data_count_cp_1(hGCZylpOryFfZNhxLZOH),
		.empty_sp_0		(qUkWgSUxlHDGwaShnpJD),
		.empty_mp_0		(AKnQHFnRxMsayGvtbpFT),
		.empty_cp_0		(EdvpzeTpOWEloDTnpLTm),
		.empty_sp_1		(vWFpyuXCRPPETqWnXLgO),
		.empty_mp_1		(dbsLvjpjMhdBsPiUgbjQ),
		.empty_cp_1		(oXZLEogkFzslyJXIZmAm),
		.dout_sp_0		(iGrqtIPPBFPUhGunhSdw),
		.dout_mp_0		(CZceBwenUmhgWecdrVuw),
		.dout_cp_0		(FODhltaveISdQIJPBJhJ),
		.dout_sp_1		(mBUfUweOiYOTkxaNfvqZ),
		.dout_mp_1		(XCEBnusbPkduEdkiHxFK),
		.dout_cp_1		(UKLUuuVquDsMMMMhkoJV),
		.rd_en_sp_0		(GVEVAzxUWjnkLWGcHbCC),
        .rd_en_mp_0     (ZOkiujEkXjtpgkcONTax),
        .rd_en_cp_0     (QcQmUnoklSTURFcjjsxj),
        .rd_en_sp_1     (artgRMUHHAMMXysfVQxf),
        .rd_en_mp_1     (CcBPKbMCVTPpuzcHaNNl),
        .rd_en_cp_1     (MQgLtHVUbOxalviVAmNV)
	);
endmodule
